
module regist_8bit_125 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]), 
        .QN() );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_124 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_123 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV4 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_83 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_82 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV1 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_83 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV4 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV4 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV4 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_82 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_81 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_122 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_80 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_81 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module cell_3_1049 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n1, n2, n3;

  LVT_XOR2HSV0 U1 ( .A1(n1), .A2(n2), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n3), .A2(t_i_1_in), .Z(n2) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n3) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n1) );
endmodule


module cell_4_146 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n2, n3, n4;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(n2) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n3) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n1) );
  LVT_XOR2HSV0 U1 ( .A1(n1), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n4) );
endmodule


module cell_4_145 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_144 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV2 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_143 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV2 U1 ( .A1(n5), .A2(n2), .A3(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_142 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_141 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10;

  LVT_INAND2HSV0 U1 ( .A1(n9), .B1(n8), .ZN(n7) );
  LVT_CLKNAND2HSV1 U2 ( .A1(n9), .A2(n5), .ZN(n6) );
  LVT_CLKNAND2HSV1 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKNHSV2 U4 ( .I(n8), .ZN(n5) );
  LVT_XNOR2HSV4 U5 ( .A1(n1), .A2(n10), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U6 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n1) );
  LVT_NAND2HSV2 U7 ( .A1(n6), .A2(n7), .ZN(n10) );
  LVT_NAND2HSV0 U8 ( .A1(b_in), .A2(a_in), .ZN(n9) );
endmodule


module cell_4_140 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  LVT_CLKNAND2HSV2 U1 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n8), .A2(n14), .ZN(n11) );
  LVT_CLKNAND2HSV2 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n13) );
  LVT_XNOR2HSV1 U4 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n12) );
  LVT_NAND2HSV2 U5 ( .A1(b_in), .A2(a_in), .ZN(n14) );
  LVT_INHSV2 U6 ( .I(n12), .ZN(n1) );
  LVT_NAND2HSV4 U7 ( .A1(n10), .A2(n11), .ZN(n15) );
  LVT_CLKNHSV2 U8 ( .I(n13), .ZN(n8) );
  LVT_NAND2HSV1 U9 ( .A1(n12), .A2(n15), .ZN(n6) );
  LVT_NAND2HSV4 U10 ( .A1(n5), .A2(n1), .ZN(n7) );
  LVT_INHSV4SR U11 ( .I(n15), .ZN(n5) );
  LVT_NAND2HSV0P5 U12 ( .A1(n13), .A2(n9), .ZN(n10) );
  LVT_INHSV0SR U13 ( .I(n14), .ZN(n9) );
endmodule


module row_1_20 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_3_1049 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_146 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(
        t_i_1_out[1]) );
  cell_4_145 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_144 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(
        t_i_1_out[3]) );
  cell_4_143 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(
        t_i_1_out[4]) );
  cell_4_142 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(
        t_i_1_out[5]) );
  cell_4_141 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_140 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_CLKNHSV1 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_146 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n1, n2;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n1) );
  LVT_XOR2HSV0 U1 ( .A1(n2), .A2(n1), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_3_1048 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1047 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1046 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1045 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1044 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV2 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_1043 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1042 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV2 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV3SR U4 ( .I(n9), .ZN(n2) );
  LVT_INHSV3 U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV4 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV4 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_146 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_146 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_1048 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1047 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1046 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1045 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1044 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1043 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1042 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_145 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_1041 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1040 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1039 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1038 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1037 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1036 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .Z(n3) );
  LVT_XOR2HSV2 U3 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n3), .A2(t_i_1_in), .ZN(n4) );
endmodule


module cell_3_1035 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_OAI21HSV2 U1 ( .A1(n6), .A2(n4), .B(n2), .ZN(t_i_out) );
  LVT_NAND2HSV4 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_NAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(n6), .ZN(n2) );
  LVT_XNOR2HSV4 U5 ( .A1(t_i_1_in), .A2(n5), .ZN(n4) );
endmodule


module row_other_145 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_145 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_1041 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1040 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1039 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1038 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1037 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1036 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1035 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_144 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_1034 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1033 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1032 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1031 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1030 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1029 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV1 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_1028 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_INHSV2 U1 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV0 U2 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV1 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2 U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV4 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_144 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_144 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_1034 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1033 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1032 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1031 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1030 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1029 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1028 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
  LVT_INHSV1SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2SR U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_143 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_1027 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1026 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1025 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1024 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1023 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1022 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1021 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_NAND2HSV0 U1 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U3 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_NAND2HSV4 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module row_other_143 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_143 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_1027 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1026 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1025 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1024 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1023 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1022 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1021 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_142 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n3), .A2(n4), .Z(t_i_out) );
endmodule


module cell_3_1020 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1019 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1018 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1017 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1016 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1015 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_1014 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9, n10;

  LVT_NAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_CLKNAND2HSV2 U3 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n9) );
  LVT_INHSV2 U5 ( .I(n8), .ZN(n5) );
  LVT_INHSV4SR U6 ( .I(n2), .ZN(n4) );
  LVT_NAND2HSV0P5 U7 ( .A1(n8), .A2(n10), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(n9), .A2(t_i_1_in), .ZN(n8) );
  LVT_NAND2HSV4 U9 ( .A1(n4), .A2(n5), .ZN(n7) );
endmodule


module row_other_142 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_142 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_1020 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1019 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1018 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1017 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1016 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1015 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1014 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_141 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4, n5, n6;

  LVT_OAI21HSV2 U1 ( .A1(n3), .A2(n5), .B(n4), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(n3), .A2(n5), .ZN(n4) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_INHSV0SR U4 ( .I(n6), .ZN(n3) );
  LVT_NAND2HSV2 U5 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_3_1013 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1012 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_1011 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1010 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_1009 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1008 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1007 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_NAND2HSV0 U1 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U3 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_NAND2HSV4 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module row_other_141 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_141 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_1013 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1012 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1011 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1010 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1009 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1008 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1007 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_140 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_1006 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_INHSV1 U5 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0P5 U6 ( .A1(n4), .A2(n7), .ZN(n5) );
endmodule


module cell_3_1005 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_1004 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1003 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_1002 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_1001 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1000 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_140 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_140 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_1006 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1005 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1004 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1003 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1002 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1001 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1000 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_20 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_20 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(
        t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), 
        .t_i_1_out(t0), .t_i_2_out(t_i_2_out[6]) );
  row_other_146 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_145 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_144 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_143 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_142 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_141 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_140 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_121 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_120 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_7bit_80 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
endmodule


module PE_20 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, 
        t_i_2_in, a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro
 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1, n1,
         n3, n4, n5, net27364, net31127, net31319, net31318, n2, n6, n7, n8,
         n9, n10;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  LVT_AO22HSV0 U11 ( .A1(mux_bq[7]), .A2(net27364), .B1(b_out[7]), .B2(
        net31127), .Z(mux_b[7]) );
  LVT_AO22HSV0 U12 ( .A1(mux_bq[6]), .A2(net27364), .B1(b_out[6]), .B2(
        net31127), .Z(mux_b[6]) );
  LVT_AO22HSV0 U13 ( .A1(mux_bq[5]), .A2(net27364), .B1(b_out[5]), .B2(
        net31127), .Z(mux_b[5]) );
  LVT_AO22HSV0 U14 ( .A1(mux_bq[4]), .A2(net27364), .B1(b_out[4]), .B2(
        net31127), .Z(mux_b[4]) );
  LVT_AO22HSV0 U15 ( .A1(mux_bq[3]), .A2(net27364), .B1(b_out[3]), .B2(
        net31127), .Z(mux_b[3]) );
  LVT_AO22HSV0 U16 ( .A1(mux_bq[2]), .A2(net27364), .B1(b_out[2]), .B2(
        net31127), .Z(mux_b[2]) );
  LVT_AO22HSV0 U17 ( .A1(mux_bq[1]), .A2(net27364), .B1(b_out[1]), .B2(
        net31127), .Z(mux_b[1]) );
  LVT_AO22HSV0 U18 ( .A1(mux_bq[0]), .A2(net27364), .B1(b_out[0]), .B2(
        net31127), .Z(mux_b[0]) );
  regist_8bit_125 u0 ( .clk(clk), .rstn(n9), .in(a_in), .out(l_a) );
  regist_8bit_124 u1 ( .clk(clk), .rstn(n9), .in(b_in), .out(b_out) );
  regist_8bit_123 u2 ( .clk(clk), .rstn(n9), .in(g_in), .out(l_g) );
  regist_1bit_83 u3 ( .clk(clk), .rstn(n9), .in(ctr), .out(l_ctr) );
  regist_1bit_82 u4 ( .clk(clk), .rstn(n9), .in(net27364), .out(ctro) );
  regist_7bit_83 u5 ( .clk(clk), .rstn(n9), .in(t_i_1_in), .out(l_t_i_1_in) );
  regist_7bit_82 u6 ( .clk(clk), .rstn(n9), .in(t_i_2_in), .out(l_t_i_2_in) );
  regist_1bit_81 u7 ( .clk(clk), .rstn(n9), .in(t_i_1_in_0), .out(l_t_i_1_in_0) );
  regist_8bit_122 u9 ( .clk(clk), .rstn(n9), .in(mux_b), .out(mux_bq) );
  regist_1bit_80 u10 ( .clk(clk), .rstn(n9), .in(net31319), .out(ti_1) );
  regist_7bit_81 u11 ( .clk(clk), .rstn(n9), .in(to_7), .out(ti_7) );
  PE_core_20 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out(t_i_2_out), .t_i_1_out_0(t_i_1_out_0)
         );
  regist_8bit_121 u12 ( .clk(clk), .rstn(n9), .in(ao), .out(a_out) );
  regist_8bit_120 u13 ( .clk(clk), .rstn(n9), .in(go), .out(g_out) );
  regist_7bit_80 u14 ( .clk(clk), .rstn(n9), .in(to), .out(t_i_1_out) );
  LVT_INHSV6 U2 ( .I(n8), .ZN(to_1) );
  LVT_INHSV0SR U3 ( .I(to_1), .ZN(net31318) );
  LVT_INHSV0SR U4 ( .I(l_ctr), .ZN(n3) );
  LVT_NAND2HSV2 U5 ( .A1(ti_7[0]), .A2(ctro), .ZN(n2) );
  LVT_CLKNAND2HSV3 U6 ( .A1(t_i_2_out[0]), .A2(n1), .ZN(n6) );
  LVT_NAND2HSV4 U7 ( .A1(n2), .A2(n6), .ZN(to_7[0]) );
  LVT_INHSV2 U8 ( .I(ctro), .ZN(n1) );
  LVT_INHSV0SR U9 ( .I(l_t_i_1_in_0), .ZN(n7) );
  LVT_NOR2HSV2 U10 ( .A1(n3), .A2(n7), .ZN(c_t_i_1_in_0) );
  LVT_INHSV6 U19 ( .I(n10), .ZN(n9) );
  LVT_MUX2NHSV4 U20 ( .I0(l_t_i_1_in_0), .I1(ti_1), .S(l_ctr), .ZN(n8) );
  LVT_INHSV2 U21 ( .I(net31318), .ZN(net31319) );
  LVT_AOI21HSV2 U22 ( .A1(n4), .A2(n5), .B(n3), .ZN(\c_t_i_1_in[0] ) );
  LVT_BUFHSV2RT U23 ( .I(n3), .Z(net31127) );
  LVT_NOR3HSV2 U24 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), .ZN(n4) );
  LVT_NOR4HSV12 U25 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(
        l_t_i_1_in[4]), .A4(l_t_i_1_in[3]), .ZN(n5) );
  LVT_INHSV2 U26 ( .I(net31127), .ZN(net27364) );
  LVT_AO22HSV4 U27 ( .A1(ti_7[2]), .A2(ctro), .B1(t_i_2_out[2]), .B2(n1), .Z(
        to_7[2]) );
  LVT_AO22HSV4 U28 ( .A1(ti_7[4]), .A2(ctro), .B1(t_i_2_out[4]), .B2(n1), .Z(
        to_7[4]) );
  LVT_AO22HSV4 U29 ( .A1(ti_7[1]), .A2(ctro), .B1(t_i_2_out[1]), .B2(n1), .Z(
        to_7[1]) );
  LVT_AO22HSV4 U30 ( .A1(ti_7[3]), .A2(ctro), .B1(t_i_2_out[3]), .B2(n1), .Z(
        to_7[3]) );
  LVT_AO22HSV4 U31 ( .A1(ti_7[5]), .A2(ctro), .B1(t_i_2_out[5]), .B2(n1), .Z(
        to_7[5]) );
  LVT_AO22HSV4 U32 ( .A1(ti_7[6]), .A2(ctro), .B1(t_i_2_out[6]), .B2(n1), .Z(
        to_7[6]) );
  LVT_INHSV2 U33 ( .I(rstn), .ZN(n10) );
endmodule


module regist_8bit_119 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_118 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_117 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_79 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_78 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV1 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_79 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV4 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV4 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV4 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV4 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_78 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
endmodule


module regist_1bit_77 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_116 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_76 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_77 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module cell_3_999 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_139 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_XOR2HSV4 U2 ( .A1(t_i_1_in), .A2(t_i_2_in), .Z(n8) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV2 U5 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_138 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_137 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_136 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n3, n4;

  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n4) );
  LVT_XNOR3HSV2 U1 ( .A1(n4), .A2(n3), .A3(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .Z(n2) );
endmodule


module cell_4_135 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10;

  LVT_INAND2HSV0 U1 ( .A1(n9), .B1(n8), .ZN(n7) );
  LVT_XNOR2HSV1 U2 ( .A1(n10), .A2(n1), .ZN(t_i_out) );
  LVT_CLKNHSV0 U3 ( .I(n8), .ZN(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_NAND2HSV2 U5 ( .A1(b_in), .A2(a_in), .ZN(n9) );
  LVT_XNOR2HSV1 U6 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n1) );
  LVT_NAND2HSV0P5 U7 ( .A1(n9), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U8 ( .A1(n6), .A2(n7), .ZN(n10) );
endmodule


module cell_4_134 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKXOR2HSV4 U2 ( .A1(n7), .A2(n8), .Z(t_i_out) );
  LVT_XOR2HSV4 U3 ( .A1(n5), .A2(n6), .Z(n7) );
endmodule


module cell_4_133 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10, n11;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n10) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n9), .A2(n10), .Z(n11) );
  LVT_XNOR2HSV1 U3 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n8) );
  LVT_INHSV2 U5 ( .I(n11), .ZN(n1) );
  LVT_NAND2HSV4 U6 ( .A1(n1), .A2(n5), .ZN(n7) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_CLKNAND2HSV1 U8 ( .A1(n11), .A2(n8), .ZN(n6) );
  LVT_INHSV2SR U9 ( .I(n8), .ZN(n5) );
endmodule


module row_1_19 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_3_999 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_139 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(
        t_i_1_out[1]) );
  cell_4_138 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_137 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(t_i_1_out[3])
         );
  cell_4_136 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(
        t_i_1_out[4]) );
  cell_4_135 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(
        t_i_1_out[5]) );
  cell_4_134 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_133 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_139 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_998 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_997 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_996 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_995 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4, n5, n6, n7;

  LVT_XNOR2HSV1 U1 ( .A1(n7), .A2(n6), .ZN(t_i_out) );
  LVT_INAND2HSV2 U2 ( .A1(n5), .B1(n2), .ZN(n4) );
  LVT_NAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n7) );
  LVT_NAND2HSV0 U5 ( .A1(n5), .A2(t_i_1_in), .ZN(n3) );
  LVT_CLKNHSV0P5 U6 ( .I(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV2 U7 ( .A1(n3), .A2(n4), .ZN(n6) );
endmodule


module cell_3_994 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_993 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_992 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  LVT_NAND2HSV2 U1 ( .A1(n9), .A2(n13), .ZN(n12) );
  LVT_INHSV2SR U2 ( .I(n14), .ZN(n6) );
  LVT_INHSV2SR U3 ( .I(n15), .ZN(n5) );
  LVT_NAND2HSV2 U4 ( .A1(n7), .A2(n8), .ZN(t_i_out) );
  LVT_NAND2HSV2 U5 ( .A1(n5), .A2(n4), .ZN(n8) );
  LVT_CLKNAND2HSV1 U6 ( .A1(n6), .A2(n15), .ZN(n7) );
  LVT_NAND2HSV0P5 U7 ( .A1(n11), .A2(n12), .ZN(n4) );
  LVT_NAND2HSV2 U8 ( .A1(n11), .A2(n12), .ZN(n14) );
  LVT_CLKNAND2HSV0 U9 ( .A1(n10), .A2(t_i_1_in), .ZN(n11) );
  LVT_NAND2HSV4 U10 ( .A1(t_m_1_in), .A2(g_in), .ZN(n15) );
  LVT_CLKNHSV2P5 U11 ( .I(t_i_1_in), .ZN(n9) );
  LVT_INHSV0SR U12 ( .I(n13), .ZN(n10) );
  LVT_NAND2HSV2 U13 ( .A1(b_in), .A2(a_in), .ZN(n13) );
endmodule


module row_other_139 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_139 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_998 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_997 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_996 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_995 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_994 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_993 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_992 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV0P5SR U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_138 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_991 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_990 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_989 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_988 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_987 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_XNOR2HSV1 U1 ( .A1(t_i_1_in), .A2(n3), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKAND2HSV2 U4 ( .A1(b_in), .A2(a_in), .Z(n3) );
endmodule


module cell_3_986 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4;

  LVT_XNOR2HSV1 U1 ( .A1(n4), .A2(n3), .ZN(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U3 ( .A1(t_i_1_in), .A2(n2), .Z(n3) );
  LVT_CLKAND2HSV2 U4 ( .A1(b_in), .A2(a_in), .Z(n2) );
endmodule


module cell_3_985 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_INAND2HSV4 U1 ( .A1(n8), .B1(n2), .ZN(n5) );
  LVT_CLKNAND2HSV3 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_INHSV4SR U4 ( .I(n6), .ZN(n2) );
  LVT_NAND2HSV1 U5 ( .A1(n8), .A2(n6), .ZN(n4) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n4), .A2(n5), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U7 ( .A1(n7), .A2(t_i_1_in), .ZN(n6) );
endmodule


module row_other_138 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_138 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_991 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_990 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_989 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_988 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_987 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_986 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_985 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_137 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_984 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_983 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_982 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_981 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_980 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_979 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_978 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV2 U2 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV0P5 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV3 U5 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV2 U6 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV4 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_137 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_137 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_984 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_983 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_982 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_981 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_980 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_979 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_978 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
  LVT_INHSV0P5SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2SR U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_136 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_977 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_976 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_975 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_974 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_973 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_972 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV0P5 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNHSV2 U4 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U5 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNHSV0 U6 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV2 U7 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U8 ( .A1(n9), .A2(n7), .ZN(n5) );
endmodule


module cell_3_971 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module row_other_136 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_136 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_977 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_976 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_975 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_974 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_973 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_972 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_971 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_135 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_970 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_969 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_968 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_967 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_966 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_965 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV1 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_964 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4;

  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n4) );
  LVT_XNOR2HSV1 U2 ( .A1(n2), .A2(t_i_1_in), .ZN(n3) );
  LVT_NAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .ZN(n2) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(n3), .ZN(t_i_out) );
endmodule


module row_other_135 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_135 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_970 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_969 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_968 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_967 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_966 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_965 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_964 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_134 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_963 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_962 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_961 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKXOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_960 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV2 U1 ( .I(n9), .ZN(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_INHSV0P5SR U5 ( .I(n10), .ZN(n4) );
  LVT_NAND2HSV2 U6 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U7 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U8 ( .A1(n4), .A2(n9), .ZN(n7) );
endmodule


module cell_3_959 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_958 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_957 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNHSV1 U1 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U4 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U5 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV0P5 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_XNOR2HSV2 U7 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_INHSV2 U8 ( .I(n7), .ZN(n4) );
endmodule


module row_other_134 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_134 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_963 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_962 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_961 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_960 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_959 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_958 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_957 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_133 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_956 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_OAI21HSV2 U1 ( .A1(t_i_1_in), .A2(n5), .B(n2), .ZN(n4) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_NAND2HSV2 U4 ( .A1(n5), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV1 U5 ( .A1(n6), .A2(n4), .ZN(t_i_out) );
endmodule


module cell_3_955 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_954 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_953 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .Z(n3) );
  LVT_XNOR2HSV4 U4 ( .A1(n3), .A2(t_i_1_in), .ZN(n4) );
endmodule


module cell_3_952 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_951 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_950 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_INHSV2SR U2 ( .I(n10), .ZN(n4) );
  LVT_NAND2HSV1 U4 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_CLKNHSV1 U5 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV0P5 U6 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U7 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_XOR2HSV2 U8 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
endmodule


module row_other_133 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_133 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_956 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_955 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_954 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_953 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_952 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_951 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_950 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_19 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_19 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(
        t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), 
        .t_i_1_out(t0), .t_i_2_out(t_i_2_out[6]) );
  row_other_139 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_138 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_137 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_136 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_135 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_134 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_133 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_115 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_114 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_7bit_76 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
endmodule


module PE_19 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, 
        t_i_2_in, a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro
 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  LVT_NOR3HSV0 U24 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), .ZN(n4) );
  regist_8bit_119 u0 ( .clk(clk), .rstn(n17), .in(a_in), .out(l_a) );
  regist_8bit_118 u1 ( .clk(clk), .rstn(n17), .in(b_in), .out(b_out) );
  regist_8bit_117 u2 ( .clk(clk), .rstn(n17), .in(g_in), .out(l_g) );
  regist_1bit_79 u3 ( .clk(clk), .rstn(n17), .in(ctr), .out(l_ctr) );
  regist_1bit_78 u4 ( .clk(clk), .rstn(n17), .in(n13), .out(ctro) );
  regist_7bit_79 u5 ( .clk(clk), .rstn(n17), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_7bit_78 u6 ( .clk(clk), .rstn(n17), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_77 u7 ( .clk(clk), .rstn(n17), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_8bit_116 u9 ( .clk(clk), .rstn(n17), .in(mux_b), .out(mux_bq) );
  regist_1bit_76 u10 ( .clk(clk), .rstn(n17), .in(to_1), .out(ti_1) );
  regist_7bit_77 u11 ( .clk(clk), .rstn(n17), .in(to_7), .out(ti_7) );
  PE_core_19 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, 
        to_7[6], n6, to_7[4:0]}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \c_t_i_1_in[0] }), .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(
        l_t_i_2_in), .a_out(ao), .g_out(go), .t_i_1_out(to), .t_i_2_out(
        t_i_2_out), .t_i_1_out_0(t_i_1_out_0) );
  regist_8bit_115 u12 ( .clk(clk), .rstn(n17), .in(ao), .out(a_out) );
  regist_8bit_114 u13 ( .clk(clk), .rstn(n17), .in(go), .out(g_out) );
  regist_7bit_76 u14 ( .clk(clk), .rstn(n17), .in(to), .out(t_i_1_out) );
  LVT_CLKNAND2HSV4 U2 ( .A1(n9), .A2(n10), .ZN(n6) );
  LVT_CLKNAND2HSV4 U3 ( .A1(n16), .A2(n15), .ZN(to_7[6]) );
  LVT_NOR2HSV0 U4 ( .A1(n2), .A2(n3), .ZN(c_t_i_1_in_0) );
  LVT_NAND2HSV0 U5 ( .A1(n9), .A2(n10), .ZN(to_7[5]) );
  LVT_NAND2HSV4 U6 ( .A1(t_i_2_out[5]), .A2(n1), .ZN(n10) );
  LVT_NAND2HSV8 U7 ( .A1(n7), .A2(n8), .ZN(to_7[1]) );
  LVT_CLKNAND2HSV8 U8 ( .A1(n11), .A2(n12), .ZN(to_7[0]) );
  LVT_INHSV4 U9 ( .I(l_t_i_1_in_0), .ZN(n2) );
  LVT_NAND2HSV2 U10 ( .A1(ti_7[1]), .A2(ctro), .ZN(n7) );
  LVT_NAND2HSV4 U11 ( .A1(t_i_2_out[1]), .A2(n1), .ZN(n8) );
  LVT_INHSV2 U12 ( .I(ctro), .ZN(n1) );
  LVT_CLKNAND2HSV1 U13 ( .A1(ti_7[5]), .A2(ctro), .ZN(n9) );
  LVT_NAND2HSV4 U14 ( .A1(ti_7[0]), .A2(ctro), .ZN(n11) );
  LVT_CLKNAND2HSV4 U15 ( .A1(t_i_2_out[0]), .A2(n1), .ZN(n12) );
  LVT_NAND2HSV2 U16 ( .A1(ti_7[6]), .A2(ctro), .ZN(n15) );
  LVT_INHSV6 U17 ( .I(n18), .ZN(n17) );
  LVT_NOR4HSV12 U18 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(
        l_t_i_1_in[4]), .A4(l_t_i_1_in[3]), .ZN(n5) );
  LVT_INHSV2 U19 ( .I(n3), .ZN(n13) );
  LVT_BUFHSV2RT U20 ( .I(n3), .Z(n14) );
  LVT_INHSV0SR U21 ( .I(l_ctr), .ZN(n3) );
  LVT_AOI21HSV2 U22 ( .A1(n4), .A2(n5), .B(n3), .ZN(\c_t_i_1_in[0] ) );
  LVT_AO22HSV2 U23 ( .A1(mux_bq[0]), .A2(n13), .B1(b_out[0]), .B2(n14), .Z(
        mux_b[0]) );
  LVT_AO22HSV2 U25 ( .A1(mux_bq[4]), .A2(n13), .B1(b_out[4]), .B2(n14), .Z(
        mux_b[4]) );
  LVT_AO22HSV2 U26 ( .A1(mux_bq[3]), .A2(l_ctr), .B1(b_out[3]), .B2(n14), .Z(
        mux_b[3]) );
  LVT_AO22HSV2 U27 ( .A1(mux_bq[1]), .A2(l_ctr), .B1(b_out[1]), .B2(n14), .Z(
        mux_b[1]) );
  LVT_AO22HSV2 U28 ( .A1(mux_bq[2]), .A2(l_ctr), .B1(b_out[2]), .B2(n14), .Z(
        mux_b[2]) );
  LVT_AO22HSV2 U29 ( .A1(mux_bq[7]), .A2(n13), .B1(b_out[7]), .B2(n14), .Z(
        mux_b[7]) );
  LVT_AO22HSV2 U30 ( .A1(mux_bq[5]), .A2(n13), .B1(b_out[5]), .B2(n14), .Z(
        mux_b[5]) );
  LVT_AO22HSV2 U31 ( .A1(mux_bq[6]), .A2(l_ctr), .B1(b_out[6]), .B2(n14), .Z(
        mux_b[6]) );
  LVT_NAND2HSV4 U32 ( .A1(t_i_2_out[6]), .A2(n1), .ZN(n16) );
  LVT_AO22HSV4 U33 ( .A1(ti_7[2]), .A2(ctro), .B1(t_i_2_out[2]), .B2(n1), .Z(
        to_7[2]) );
  LVT_AO22HSV4 U34 ( .A1(ti_7[3]), .A2(ctro), .B1(t_i_2_out[3]), .B2(n1), .Z(
        to_7[3]) );
  LVT_AO22HSV4 U35 ( .A1(ti_7[4]), .A2(ctro), .B1(t_i_2_out[4]), .B2(n1), .Z(
        to_7[4]) );
  LVT_MOAI22HSV4 U36 ( .A1(l_ctr), .A2(n2), .B1(l_ctr), .B2(ti_1), .ZN(to_1)
         );
  LVT_INHSV2 U37 ( .I(rstn), .ZN(n18) );
endmodule


module regist_8bit_113 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_112 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_111 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_75 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_74 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_75 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_74 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_73 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_110 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_72 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_73 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module cell_3_949 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_132 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_131 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV2 U1 ( .A1(n5), .A2(n2), .A3(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_130 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_129 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_128 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_127 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n5, n6, n7;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n7) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n6), .ZN(n2) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U3 ( .A1(n7), .A2(n2), .ZN(t_i_out) );
endmodule


module cell_4_126 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  LVT_INAND2HSV0 U1 ( .A1(n13), .B1(n12), .ZN(n11) );
  LVT_CLKNAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n12) );
  LVT_INHSV2 U3 ( .I(n12), .ZN(n9) );
  LVT_XNOR2HSV1 U4 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n8) );
  LVT_NAND2HSV4 U5 ( .A1(n1), .A2(n5), .ZN(n7) );
  LVT_INHSV2 U6 ( .I(n14), .ZN(n1) );
  LVT_NAND2HSV0P5 U7 ( .A1(n14), .A2(n8), .ZN(n6) );
  LVT_CLKNAND2HSV3 U8 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV3SR U9 ( .I(n8), .ZN(n5) );
  LVT_NAND2HSV0P5 U10 ( .A1(n13), .A2(n9), .ZN(n10) );
  LVT_NAND2HSV2 U11 ( .A1(n10), .A2(n11), .ZN(n14) );
  LVT_NAND2HSV0 U12 ( .A1(b_in), .A2(a_in), .ZN(n13) );
endmodule


module row_1_18 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_3_949 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_132 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(
        t_i_1_out[1]) );
  cell_4_131 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_130 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(
        t_i_1_out[3]) );
  cell_4_129 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(
        t_i_1_out[4]) );
  cell_4_128 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(
        t_i_1_out[5]) );
  cell_4_127 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_126 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
endmodule


module cell_2_132 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_948 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_947 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_946 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_945 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_944 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_943 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_INHSV2SR U5 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0P5 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_942 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV2 U4 ( .I(n7), .ZN(n4) );
  LVT_INHSV3SR U5 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV0 U6 ( .A1(n7), .A2(n9), .ZN(n5) );
  LVT_NAND2HSV4 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_132 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_132 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_948 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_947 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_946 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_945 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_944 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_943 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_942 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_131 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_941 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_940 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_939 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U5 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_938 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_937 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_936 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module cell_3_935 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2SR U4 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV1 U6 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNAND2HSV0 U7 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2SR U8 ( .I(n7), .ZN(n4) );
endmodule


module row_other_131 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_131 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_941 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_940 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_939 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_938 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_937 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_936 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_935 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_130 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_934 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_933 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_932 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_931 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_930 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_929 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_928 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U2 ( .A1(n7), .A2(n9), .ZN(n5) );
  LVT_INHSV3SR U4 ( .I(n9), .ZN(n2) );
  LVT_CLKNHSV4 U5 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_NAND2HSV4 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_130 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_130 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_934 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_933 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_932 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_931 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_930 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_929 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_928 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_129 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_927 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_926 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_925 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_XOR2HSV0 U2 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNHSV0P5 U5 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV2 U6 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U7 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV2 U8 ( .I(n8), .ZN(n4) );
endmodule


module cell_3_924 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_923 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_NAND2HSV2 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV1 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_922 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_NAND2HSV0P5 U1 ( .A1(n5), .A2(t_i_1_in), .ZN(n2) );
  LVT_OAI21HSV2 U2 ( .A1(t_i_1_in), .A2(n5), .B(n2), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XNOR2HSV4 U5 ( .A1(n6), .A2(n4), .ZN(t_i_out) );
endmodule


module cell_3_921 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV2 U1 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV4 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_NAND2HSV2 U5 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV4 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV3SR U7 ( .I(n9), .ZN(n2) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_129 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_129 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_927 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_926 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_925 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_924 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_923 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_922 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_921 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_128 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_920 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_919 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_918 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_917 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_916 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_915 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_914 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U1 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV3 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV2 U4 ( .I(n7), .ZN(n4) );
  LVT_INHSV3SR U5 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV4 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_128 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_128 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_920 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_919 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_918 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_917 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_916 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_915 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_914 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_127 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_913 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_912 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_911 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_910 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_909 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_908 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_907 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module row_other_127 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_127 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_913 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_912 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_911 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_910 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_909 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_908 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_907 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_126 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4, n5, n6, n7;

  LVT_INAND2HSV2 U1 ( .A1(n6), .B1(n7), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(n3), .A2(n6), .ZN(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(n4), .A2(n5), .ZN(t_i_out) );
  LVT_INHSV0SR U4 ( .I(n7), .ZN(n3) );
  LVT_NAND2HSV2 U5 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_NAND2HSV0P5 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_906 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n10) );
  LVT_OAI21HSV2 U1 ( .A1(n8), .A2(t_i_1_in), .B(n9), .ZN(n11) );
  LVT_NAND2HSV0P5 U2 ( .A1(n12), .A2(n5), .ZN(n6) );
  LVT_CLKNAND2HSV1 U4 ( .A1(n4), .A2(n11), .ZN(n7) );
  LVT_CLKNAND2HSV0 U5 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV0SR U6 ( .I(n12), .ZN(n4) );
  LVT_INHSV0SR U7 ( .I(n11), .ZN(n5) );
  LVT_NAND2HSV0P5 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n12) );
  LVT_NAND2HSV2 U9 ( .A1(n8), .A2(t_i_1_in), .ZN(n9) );
  LVT_INHSV2 U10 ( .I(n10), .ZN(n8) );
endmodule


module cell_3_905 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module cell_3_904 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XNOR2HSV4 U1 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV0P5 U2 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV2 U4 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV1SR U6 ( .I(n9), .ZN(n2) );
  LVT_INHSV2 U7 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV0P5 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
endmodule


module cell_3_903 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_902 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_INHSV2SR U4 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV0 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U6 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U7 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV2 U8 ( .I(n8), .ZN(n4) );
endmodule


module cell_3_901 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_900 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module row_other_126 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_126 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_906 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_905 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_904 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_903 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_902 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_901 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_900 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_18 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_18 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(
        t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), 
        .t_i_1_out(t0), .t_i_2_out(t_i_2_out[6]) );
  row_other_132 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_131 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_130 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_129 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_128 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_127 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_126 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_109 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_108 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_72 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module PE_18 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, 
        t_i_2_in, a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro
 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  LVT_NOR3HSV0 U24 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), .ZN(n14) );
  regist_8bit_113 u0 ( .clk(clk), .rstn(rstn), .in(a_in), .out(l_a) );
  regist_8bit_112 u1 ( .clk(clk), .rstn(rstn), .in(b_in), .out(b_out) );
  regist_8bit_111 u2 ( .clk(clk), .rstn(rstn), .in(g_in), .out(l_g) );
  regist_1bit_75 u3 ( .clk(clk), .rstn(rstn), .in(ctr), .out(l_ctr) );
  regist_1bit_74 u4 ( .clk(clk), .rstn(rstn), .in(n12), .out(ctro) );
  regist_7bit_75 u5 ( .clk(clk), .rstn(rstn), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_7bit_74 u6 ( .clk(clk), .rstn(rstn), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_73 u7 ( .clk(clk), .rstn(rstn), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_8bit_110 u9 ( .clk(clk), .rstn(rstn), .in(mux_b), .out(mux_bq) );
  regist_1bit_72 u10 ( .clk(clk), .rstn(rstn), .in(n6), .out(ti_1) );
  regist_7bit_73 u11 ( .clk(clk), .rstn(rstn), .in(to_7), .out(ti_7) );
  PE_core_18 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out(t_i_2_out), .t_i_1_out_0(t_i_1_out_0)
         );
  regist_8bit_109 u12 ( .clk(clk), .rstn(rstn), .in(ao), .out(a_out) );
  regist_8bit_108 u13 ( .clk(clk), .rstn(rstn), .in(go), .out(g_out) );
  regist_7bit_72 u14 ( .clk(clk), .rstn(rstn), .in(to), .out(t_i_1_out) );
  LVT_MOAI22HSV0 U2 ( .A1(l_ctr), .A2(n16), .B1(ti_1), .B2(l_ctr), .ZN(n6) );
  LVT_INHSV4SR U3 ( .I(l_t_i_1_in_0), .ZN(n16) );
  LVT_MOAI22HSV4 U4 ( .A1(l_ctr), .A2(n16), .B1(ti_1), .B2(l_ctr), .ZN(to_1)
         );
  LVT_INHSV2P5 U5 ( .I(l_ctr), .ZN(n15) );
  LVT_INHSV2 U6 ( .I(n15), .ZN(n7) );
  LVT_AOI21HSV2 U7 ( .A1(n14), .A2(n13), .B(n15), .ZN(\c_t_i_1_in[0] ) );
  LVT_NOR4HSV12 U8 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(l_t_i_1_in[4]), .A4(l_t_i_1_in[3]), .ZN(n13) );
  LVT_NAND2HSV0P5 U9 ( .A1(ti_7[0]), .A2(ctro), .ZN(n8) );
  LVT_CLKNAND2HSV3 U10 ( .A1(t_i_2_out[0]), .A2(n17), .ZN(n9) );
  LVT_NAND2HSV4 U11 ( .A1(n8), .A2(n9), .ZN(to_7[0]) );
  LVT_INHSV2 U12 ( .I(ctro), .ZN(n17) );
  LVT_CLKNAND2HSV1 U13 ( .A1(ti_7[4]), .A2(ctro), .ZN(n10) );
  LVT_CLKNAND2HSV3 U14 ( .A1(t_i_2_out[4]), .A2(n17), .ZN(n11) );
  LVT_NAND2HSV4 U15 ( .A1(n10), .A2(n11), .ZN(to_7[4]) );
  LVT_NOR2HSV0 U16 ( .A1(n16), .A2(n15), .ZN(c_t_i_1_in_0) );
  LVT_CLKNHSV1 U17 ( .I(n15), .ZN(n12) );
  LVT_AO22HSV2 U18 ( .A1(mux_bq[4]), .A2(n12), .B1(b_out[4]), .B2(n15), .Z(
        mux_b[4]) );
  LVT_AO22HSV2 U19 ( .A1(mux_bq[0]), .A2(n12), .B1(b_out[0]), .B2(n15), .Z(
        mux_b[0]) );
  LVT_AO22HSV2 U20 ( .A1(mux_bq[1]), .A2(n12), .B1(b_out[1]), .B2(n15), .Z(
        mux_b[1]) );
  LVT_AO22HSV2 U21 ( .A1(mux_bq[2]), .A2(n12), .B1(b_out[2]), .B2(n15), .Z(
        mux_b[2]) );
  LVT_AO22HSV2 U22 ( .A1(mux_bq[3]), .A2(n12), .B1(b_out[3]), .B2(n15), .Z(
        mux_b[3]) );
  LVT_AO22HSV2 U23 ( .A1(mux_bq[5]), .A2(n7), .B1(b_out[5]), .B2(n15), .Z(
        mux_b[5]) );
  LVT_AO22HSV2 U25 ( .A1(mux_bq[7]), .A2(n7), .B1(b_out[7]), .B2(n15), .Z(
        mux_b[7]) );
  LVT_AO22HSV2 U26 ( .A1(mux_bq[6]), .A2(n7), .B1(b_out[6]), .B2(n15), .Z(
        mux_b[6]) );
  LVT_AO22HSV4 U27 ( .A1(ti_7[1]), .A2(ctro), .B1(t_i_2_out[1]), .B2(n17), .Z(
        to_7[1]) );
  LVT_AO22HSV4 U28 ( .A1(ti_7[2]), .A2(ctro), .B1(t_i_2_out[2]), .B2(n17), .Z(
        to_7[2]) );
  LVT_AO22HSV4 U29 ( .A1(ti_7[3]), .A2(ctro), .B1(t_i_2_out[3]), .B2(n17), .Z(
        to_7[3]) );
  LVT_AO22HSV4 U30 ( .A1(ti_7[6]), .A2(ctro), .B1(t_i_2_out[6]), .B2(n17), .Z(
        to_7[6]) );
  LVT_AO22HSV4 U31 ( .A1(ti_7[5]), .A2(ctro), .B1(t_i_2_out[5]), .B2(n17), .Z(
        to_7[5]) );
endmodule


module regist_8bit_107 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_106 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_105 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_71 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_70 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_71 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV4 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_70 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_69 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_104 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_68 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_69 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module cell_3_899 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_CLKNAND2HSV1 U2 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_CLKNHSV0 U4 ( .I(n8), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_4_125 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV4 U3 ( .A1(t_i_1_in), .A2(t_i_2_in), .Z(n8) );
  LVT_XOR2HSV0 U5 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_124 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_123 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_122 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_121 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n2), .A3(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_120 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10, n11;

  LVT_XNOR2HSV1 U1 ( .A1(n11), .A2(n1), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .ZN(n10) );
  LVT_XNOR2HSV1 U3 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n1) );
  LVT_CLKNHSV0P5 U4 ( .I(n9), .ZN(n6) );
  LVT_NAND2HSV0 U5 ( .A1(n5), .A2(n9), .ZN(n8) );
  LVT_CLKNAND2HSV1 U6 ( .A1(n10), .A2(n6), .ZN(n7) );
  LVT_NAND2HSV2 U7 ( .A1(n7), .A2(n8), .ZN(n11) );
  LVT_INHSV0SR U8 ( .I(n10), .ZN(n5) );
  LVT_NAND2HSV0P5 U9 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
endmodule


module cell_4_119 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10, n11;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n10) );
  LVT_INHSV2SR U1 ( .I(n11), .ZN(n5) );
  LVT_NAND2HSV2 U2 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_NAND2HSV2 U3 ( .A1(n1), .A2(n5), .ZN(n7) );
  LVT_CLKNAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV1 U6 ( .A1(n8), .A2(n11), .ZN(n6) );
  LVT_XOR2HSV4 U7 ( .A1(n9), .A2(n10), .Z(n11) );
  LVT_INHSV2 U8 ( .I(n8), .ZN(n1) );
  LVT_XNOR2HSV1 U9 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n8) );
endmodule


module row_1_17 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_3_899 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_125 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(
        t_i_1_out[1]) );
  cell_4_124 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_123 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(
        t_i_1_out[3]) );
  cell_4_122 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(
        t_i_1_out[4]) );
  cell_4_121 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(
        t_i_1_out[5]) );
  cell_4_120 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_119 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_125 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_898 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_897 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_896 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_895 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_894 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_893 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_892 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module row_other_125 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_125 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_898 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_897 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_896 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_895 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_894 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_893 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_892 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_124 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_891 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_890 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_889 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_888 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_887 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_886 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_885 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV3SR U1 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV3 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNHSV2P5 U5 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_CLKNAND2HSV1 U7 ( .A1(n7), .A2(n9), .ZN(n5) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_124 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_124 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_891 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_890 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_889 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_888 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_887 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_886 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_885 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_123 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_884 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV1 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_883 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_882 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_881 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_880 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_879 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_878 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_123 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_123 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_884 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_883 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_882 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_881 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_880 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_879 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_878 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_122 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_877 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_876 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(g_in), .A2(t_m_1_in), .ZN(n6) );
endmodule


module cell_3_875 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_874 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_873 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(g_in), .A2(t_m_1_in), .ZN(n6) );
endmodule


module cell_3_872 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_871 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV2SR U1 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV0 U2 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV2 U4 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV4 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV1 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_122 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_122 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_877 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_876 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_875 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_874 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_873 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_872 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_871 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_121 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4, n5, n6, n7, n8;

  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n7) );
  LVT_NAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV0P5SR U3 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(n8), .A2(n4), .ZN(n5) );
  LVT_CLKNAND2HSV0 U5 ( .A1(n3), .A2(n7), .ZN(n6) );
  LVT_NAND2HSV2 U6 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV0SR U7 ( .I(n8), .ZN(n3) );
endmodule


module cell_3_870 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_869 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_868 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_867 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_866 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_865 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_864 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module row_other_121 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_121 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_870 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_869 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_868 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_867 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_866 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_865 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_864 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_120 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_863 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_862 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_861 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_OAI21HSV2 U1 ( .A1(t_i_1_in), .A2(n5), .B(n2), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(n5), .A2(t_i_1_in), .ZN(n2) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XNOR2HSV4 U5 ( .A1(n6), .A2(n4), .ZN(t_i_out) );
endmodule


module cell_3_860 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_859 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_858 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_XOR2HSV2 U5 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_INHSV2 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_857 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNHSV2 U4 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNHSV2 U6 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV1 U7 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_120 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_120 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_863 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_862 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_861 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_860 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_859 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_858 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_857 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_119 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_856 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_855 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_854 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_853 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_852 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_851 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_850 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module row_other_119 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_119 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_856 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_855 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_854 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_853 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_852 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_851 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_850 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_17 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_17 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(
        t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), 
        .t_i_1_out(t0), .t_i_2_out(t_i_2_out[6]) );
  row_other_125 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_124 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_123 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_122 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_121 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_120 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_119 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_103 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_102 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_68 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module PE_17 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, 
        t_i_2_in, a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro
 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   n22, l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1,
         n6, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  regist_8bit_107 u0 ( .clk(clk), .rstn(rstn), .in(a_in), .out(l_a) );
  regist_8bit_106 u1 ( .clk(clk), .rstn(rstn), .in(b_in), .out(b_out) );
  regist_8bit_105 u2 ( .clk(clk), .rstn(rstn), .in(g_in), .out(l_g) );
  regist_1bit_71 u3 ( .clk(clk), .rstn(rstn), .in(ctr), .out(l_ctr) );
  regist_1bit_70 u4 ( .clk(clk), .rstn(rstn), .in(n14), .out(ctro) );
  regist_7bit_71 u5 ( .clk(clk), .rstn(rstn), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_7bit_70 u6 ( .clk(clk), .rstn(rstn), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_69 u7 ( .clk(clk), .rstn(rstn), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_8bit_104 u9 ( .clk(clk), .rstn(rstn), .in(mux_b), .out(mux_bq) );
  regist_1bit_68 u10 ( .clk(clk), .rstn(rstn), .in(n13), .out(ti_1) );
  regist_7bit_69 u11 ( .clk(clk), .rstn(rstn), .in(to_7), .out(ti_7) );
  PE_core_17 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out({t_i_2_out[6:1], n22}), .t_i_1_out_0(
        t_i_1_out_0) );
  regist_8bit_103 u12 ( .clk(clk), .rstn(rstn), .in(ao), .out(a_out) );
  regist_8bit_102 u13 ( .clk(clk), .rstn(rstn), .in(go), .out(g_out) );
  regist_7bit_68 u14 ( .clk(clk), .rstn(rstn), .in(to), .out(t_i_1_out) );
  LVT_NAND2HSV4 U2 ( .A1(t_i_2_out[1]), .A2(n21), .ZN(n16) );
  LVT_AOI21HSV1 U3 ( .A1(n18), .A2(n17), .B(n19), .ZN(\c_t_i_1_in[0] ) );
  LVT_AO22HSV1 U4 ( .A1(mux_bq[7]), .A2(n14), .B1(b_out[7]), .B2(n19), .Z(
        mux_b[7]) );
  LVT_AO22HSV1 U5 ( .A1(mux_bq[6]), .A2(n14), .B1(b_out[6]), .B2(n19), .Z(
        mux_b[6]) );
  LVT_INHSV0SR U6 ( .I(n22), .ZN(n6) );
  LVT_INHSV2 U7 ( .I(n6), .ZN(t_i_2_out[0]) );
  LVT_NOR2HSV0 U8 ( .A1(n20), .A2(n19), .ZN(c_t_i_1_in_0) );
  LVT_NOR3HSV2 U9 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), 
        .ZN(n18) );
  LVT_CLKNAND2HSV8 U10 ( .A1(n16), .A2(n15), .ZN(to_7[1]) );
  LVT_INHSV4 U11 ( .I(l_t_i_1_in_0), .ZN(n20) );
  LVT_NAND2HSV8 U12 ( .A1(n10), .A2(n11), .ZN(to_7[0]) );
  LVT_NOR4HSV12 U13 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(
        l_t_i_1_in[4]), .A4(l_t_i_1_in[3]), .ZN(n17) );
  LVT_INHSV2 U14 ( .I(ctro), .ZN(n21) );
  LVT_NAND2HSV2 U15 ( .A1(ti_7[0]), .A2(ctro), .ZN(n10) );
  LVT_NAND2HSV2 U16 ( .A1(ti_7[6]), .A2(ctro), .ZN(n8) );
  LVT_NAND2HSV2 U17 ( .A1(t_i_2_out[6]), .A2(n21), .ZN(n9) );
  LVT_NAND2HSV4 U18 ( .A1(n8), .A2(n9), .ZN(to_7[6]) );
  LVT_CLKNAND2HSV4 U19 ( .A1(n22), .A2(n21), .ZN(n11) );
  LVT_AO22HSV1 U20 ( .A1(mux_bq[0]), .A2(n14), .B1(b_out[0]), .B2(n19), .Z(
        mux_b[0]) );
  LVT_AO22HSV1 U21 ( .A1(mux_bq[1]), .A2(n14), .B1(b_out[1]), .B2(n19), .Z(
        mux_b[1]) );
  LVT_AO22HSV1 U22 ( .A1(mux_bq[2]), .A2(n14), .B1(b_out[2]), .B2(n19), .Z(
        mux_b[2]) );
  LVT_AO22HSV1 U23 ( .A1(mux_bq[3]), .A2(n14), .B1(b_out[3]), .B2(n19), .Z(
        mux_b[3]) );
  LVT_AO22HSV1 U24 ( .A1(mux_bq[4]), .A2(n14), .B1(b_out[4]), .B2(n19), .Z(
        mux_b[4]) );
  LVT_AO22HSV0 U25 ( .A1(mux_bq[5]), .A2(n14), .B1(b_out[5]), .B2(n19), .Z(
        mux_b[5]) );
  LVT_INHSV0SR U26 ( .I(to_1), .ZN(n12) );
  LVT_INHSV2 U27 ( .I(n12), .ZN(n13) );
  LVT_INHSV0P5 U28 ( .I(l_ctr), .ZN(n19) );
  LVT_INHSV0SR U29 ( .I(n19), .ZN(n14) );
  LVT_NAND2HSV2 U30 ( .A1(ti_7[1]), .A2(ctro), .ZN(n15) );
  LVT_AO22HSV4 U31 ( .A1(ti_7[2]), .A2(ctro), .B1(t_i_2_out[2]), .B2(n21), .Z(
        to_7[2]) );
  LVT_AO22HSV4 U32 ( .A1(ti_7[3]), .A2(ctro), .B1(t_i_2_out[3]), .B2(n21), .Z(
        to_7[3]) );
  LVT_AO22HSV4 U33 ( .A1(ti_7[4]), .A2(ctro), .B1(t_i_2_out[4]), .B2(n21), .Z(
        to_7[4]) );
  LVT_AO22HSV4 U34 ( .A1(ti_7[5]), .A2(ctro), .B1(t_i_2_out[5]), .B2(n21), .Z(
        to_7[5]) );
  LVT_MOAI22HSV4 U35 ( .A1(l_ctr), .A2(n20), .B1(l_ctr), .B2(ti_1), .ZN(to_1)
         );
endmodule


module regist_8bit_101 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_100 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_99 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_67 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_66 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV1 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_67 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_66 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
endmodule


module regist_1bit_65 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_98 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_64 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_65 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module cell_3_849 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_118 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV2 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_NAND2HSV2 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_117 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_116 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_115 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n7), .A2(n8), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_114 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n3, n5, n6, n7, n8, n9, n10;

  LVT_XNOR2HSV2 U1 ( .A1(n7), .A2(n10), .ZN(t_i_out) );
  LVT_INHSV0P5 U2 ( .I(n9), .ZN(n3) );
  LVT_NAND2HSV0 U3 ( .A1(n8), .A2(n9), .ZN(n5) );
  LVT_CLKNAND2HSV1 U4 ( .A1(n1), .A2(n3), .ZN(n6) );
  LVT_NAND2HSV2 U5 ( .A1(n5), .A2(n6), .ZN(n10) );
  LVT_INHSV0 U6 ( .I(n8), .ZN(n1) );
  LVT_CLKAND2HSV2 U7 ( .A1(b_in), .A2(a_in), .Z(n8) );
  LVT_NAND2HSV0P5 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV1 U9 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n7) );
endmodule


module cell_4_113 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n5, n6, n7;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n7) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n6), .ZN(n2) );
  LVT_XNOR2HSV4 U2 ( .A1(n7), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_112 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n12) );
  LVT_CLKNAND2HSV2 U2 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INAND2HSV0 U3 ( .A1(n13), .B1(n12), .ZN(n11) );
  LVT_NAND2HSV2 U4 ( .A1(n10), .A2(n11), .ZN(n14) );
  LVT_NAND2HSV2 U5 ( .A1(n9), .A2(n13), .ZN(n10) );
  LVT_INHSV2 U6 ( .I(n14), .ZN(n1) );
  LVT_XNOR2HSV1 U7 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n8) );
  LVT_CLKNHSV2 U8 ( .I(n12), .ZN(n9) );
  LVT_NAND2HSV1 U9 ( .A1(n14), .A2(n8), .ZN(n6) );
  LVT_CLKNAND2HSV3 U10 ( .A1(n1), .A2(n5), .ZN(n7) );
  LVT_CLKNHSV2 U11 ( .I(n8), .ZN(n5) );
  LVT_NAND2HSV0 U12 ( .A1(b_in), .A2(a_in), .ZN(n13) );
endmodule


module row_1_16 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_3_849 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_118 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(t_i_1_out[1])
         );
  cell_4_117 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_116 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(
        t_i_1_out[3]) );
  cell_4_115 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(
        t_i_1_out[4]) );
  cell_4_114 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(
        t_i_1_out[5]) );
  cell_4_113 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_112 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
  LVT_CLKNHSV2 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_118 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_848 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_847 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_846 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_845 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_844 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_XNOR2HSV1 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_843 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4, n5, n6, n7, n8;

  LVT_NAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U2 ( .A1(n6), .A2(n3), .ZN(n4) );
  LVT_NAND2HSV2 U3 ( .A1(n2), .A2(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(n5), .ZN(n7) );
  LVT_INHSV2 U5 ( .I(n6), .ZN(n2) );
  LVT_INHSV2 U6 ( .I(t_i_1_in), .ZN(n3) );
  LVT_CLKAND2HSV2 U7 ( .A1(b_in), .A2(a_in), .Z(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(n7), .ZN(t_i_out) );
endmodule


module cell_3_842 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U2 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U5 ( .I(n9), .ZN(n2) );
  LVT_INHSV2 U6 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV1 U7 ( .A1(n7), .A2(n9), .ZN(n5) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_118 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_118 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_848 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_847 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_846 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_845 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_844 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_843 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_842 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_117 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_841 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_840 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_839 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_838 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_837 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_836 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_835 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_117 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_117 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_841 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_840 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_839 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_838 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_837 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_836 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_835 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_116 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_834 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_833 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_832 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_831 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_830 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_829 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_828 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV4 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module row_other_116 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_116 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_834 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_833 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_832 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_831 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_830 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_829 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_828 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV0SR U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_115 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_827 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_826 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_825 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_824 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_823 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_822 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_821 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV3SR U2 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_NAND2HSV4 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV4 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_115 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_115 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_827 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_826 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_825 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_824 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_823 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_822 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_821 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_114 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_820 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_819 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_818 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_817 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV0P5 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNHSV2 U5 ( .I(n9), .ZN(n2) );
  LVT_INHSV2 U6 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV1 U7 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNAND2HSV0 U8 ( .A1(g_in), .A2(t_m_1_in), .ZN(n9) );
endmodule


module cell_3_816 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_815 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_814 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV1 U2 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV0 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV3 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV4 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_114 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_114 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_820 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_819 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_818 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_817 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_816 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_815 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_814 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_113 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_813 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_812 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U2 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
  LVT_INHSV2 U4 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV0P5 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV0P5 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV2 U7 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNHSV2 U8 ( .I(n9), .ZN(n2) );
endmodule


module cell_3_811 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKNHSV0P5 U4 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_XOR2HSV2 U6 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
endmodule


module cell_3_810 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_809 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_CLKAND2HSV2 U1 ( .A1(b_in), .A2(a_in), .Z(n3) );
  LVT_XNOR2HSV4 U2 ( .A1(n3), .A2(t_i_1_in), .ZN(n4) );
  LVT_XOR2HSV2 U3 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_808 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_807 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_OAI21HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .B(n5), .ZN(n7) );
  LVT_CLKNAND2HSV3 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U3 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_INHSV2 U5 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module row_other_113 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_113 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_813 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_812 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_811 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_810 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_809 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_808 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_807 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_112 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4, n5, n6;

  LVT_OAI21HSV2 U1 ( .A1(n3), .A2(n5), .B(n4), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U3 ( .A1(n3), .A2(n5), .ZN(n4) );
  LVT_INHSV0SR U4 ( .I(n6), .ZN(n3) );
  LVT_NAND2HSV0P5 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_806 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV2 U1 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_CLKNAND2HSV1 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_CLKNHSV0P5 U4 ( .I(n9), .ZN(n5) );
  LVT_INHSV0P5SR U5 ( .I(n10), .ZN(n4) );
  LVT_NAND2HSV0P5 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV0P5 U7 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_CLKNAND2HSV0 U8 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
endmodule


module cell_3_805 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_XNOR2HSV1 U1 ( .A1(n3), .A2(t_i_1_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKAND2HSV2 U4 ( .A1(b_in), .A2(a_in), .Z(n3) );
endmodule


module cell_3_804 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_803 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNHSV0P5 U1 ( .I(n9), .ZN(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_INHSV0SR U4 ( .I(n10), .ZN(n4) );
  LVT_NAND2HSV0P5 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV0P5 U6 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0P5 U7 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_CLKNAND2HSV0 U8 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
endmodule


module cell_3_802 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_801 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_XOR2HSV0 U2 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U6 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV2 U7 ( .I(n8), .ZN(n4) );
  LVT_INHSV2 U8 ( .I(t_i_1_in), .ZN(n5) );
endmodule


module cell_3_800 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_INHSV2 U2 ( .I(n10), .ZN(n4) );
  LVT_CLKNHSV2 U4 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV2 U5 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U6 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0P5 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_XOR2HSV2 U8 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
endmodule


module row_other_112 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_112 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_806 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_805 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_804 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_803 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_802 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_801 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_800 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_16 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_16 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(
        t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), 
        .t_i_1_out(t0), .t_i_2_out(t_i_2_out[6]) );
  row_other_118 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_117 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_116 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_115 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_114 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_113 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_112 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_97 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_96 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_7bit_64 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module PE_16 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, 
        t_i_2_in, a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro
 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  LVT_NOR3HSV0 U24 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), .ZN(n17) );
  regist_8bit_101 u0 ( .clk(clk), .rstn(n14), .in(a_in), .out(l_a) );
  regist_8bit_100 u1 ( .clk(clk), .rstn(n14), .in(b_in), .out(b_out) );
  regist_8bit_99 u2 ( .clk(clk), .rstn(n14), .in(g_in), .out(l_g) );
  regist_1bit_67 u3 ( .clk(clk), .rstn(n14), .in(ctr), .out(l_ctr) );
  regist_1bit_66 u4 ( .clk(clk), .rstn(n14), .in(n11), .out(ctro) );
  regist_7bit_67 u5 ( .clk(clk), .rstn(n14), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_7bit_66 u6 ( .clk(clk), .rstn(n14), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_65 u7 ( .clk(clk), .rstn(n14), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_8bit_98 u9 ( .clk(clk), .rstn(n14), .in(mux_b), .out(mux_bq) );
  regist_1bit_64 u10 ( .clk(clk), .rstn(n14), .in(n10), .out(ti_1) );
  regist_7bit_65 u11 ( .clk(clk), .rstn(n14), .in(to_7), .out(ti_7) );
  PE_core_16 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out(t_i_2_out), .t_i_1_out_0(t_i_1_out_0)
         );
  regist_8bit_97 u12 ( .clk(clk), .rstn(n14), .in(ao), .out(a_out) );
  regist_8bit_96 u13 ( .clk(clk), .rstn(n14), .in(go), .out(g_out) );
  regist_7bit_64 u14 ( .clk(clk), .rstn(n14), .in(to), .out(t_i_1_out) );
  LVT_NAND2HSV8 U2 ( .A1(n6), .A2(n7), .ZN(to_7[0]) );
  LVT_NOR4HSV12 U3 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(l_t_i_1_in[4]), .A4(l_t_i_1_in[3]), .ZN(n16) );
  LVT_NAND2HSV2 U4 ( .A1(ti_7[1]), .A2(ctro), .ZN(n12) );
  LVT_NAND2HSV4 U5 ( .A1(t_i_2_out[1]), .A2(n20), .ZN(n13) );
  LVT_CLKNAND2HSV4 U6 ( .A1(n8), .A2(n9), .ZN(to_7[5]) );
  LVT_NAND2HSV2 U7 ( .A1(t_i_2_out[5]), .A2(n20), .ZN(n9) );
  LVT_INHSV2 U8 ( .I(ctro), .ZN(n20) );
  LVT_NAND2HSV2 U9 ( .A1(ti_7[0]), .A2(ctro), .ZN(n6) );
  LVT_CLKNAND2HSV3 U10 ( .A1(t_i_2_out[0]), .A2(n20), .ZN(n7) );
  LVT_NAND2HSV2 U11 ( .A1(ti_7[5]), .A2(ctro), .ZN(n8) );
  LVT_INHSV6 U12 ( .I(n15), .ZN(n14) );
  LVT_INHSV2 U13 ( .I(l_ctr), .ZN(n18) );
  LVT_INHSV4SR U14 ( .I(l_t_i_1_in_0), .ZN(n19) );
  LVT_MOAI22HSV0 U15 ( .A1(n11), .A2(n19), .B1(ti_1), .B2(l_ctr), .ZN(n10) );
  LVT_NOR2HSV0 U16 ( .A1(n19), .A2(n18), .ZN(c_t_i_1_in_0) );
  LVT_INHSV2 U17 ( .I(n18), .ZN(n11) );
  LVT_AOI21HSV2 U18 ( .A1(n17), .A2(n16), .B(n18), .ZN(\c_t_i_1_in[0] ) );
  LVT_CLKNAND2HSV8 U19 ( .A1(n13), .A2(n12), .ZN(to_7[1]) );
  LVT_AO22HSV2 U20 ( .A1(mux_bq[0]), .A2(n11), .B1(b_out[0]), .B2(n18), .Z(
        mux_b[0]) );
  LVT_AO22HSV2 U21 ( .A1(mux_bq[1]), .A2(n11), .B1(b_out[1]), .B2(n18), .Z(
        mux_b[1]) );
  LVT_AO22HSV2 U22 ( .A1(mux_bq[2]), .A2(n11), .B1(b_out[2]), .B2(n18), .Z(
        mux_b[2]) );
  LVT_AO22HSV2 U23 ( .A1(mux_bq[3]), .A2(n11), .B1(b_out[3]), .B2(n18), .Z(
        mux_b[3]) );
  LVT_AO22HSV2 U25 ( .A1(mux_bq[4]), .A2(n11), .B1(b_out[4]), .B2(n18), .Z(
        mux_b[4]) );
  LVT_AO22HSV2 U26 ( .A1(mux_bq[5]), .A2(n11), .B1(b_out[5]), .B2(n18), .Z(
        mux_b[5]) );
  LVT_AO22HSV2 U27 ( .A1(mux_bq[6]), .A2(n11), .B1(b_out[6]), .B2(n18), .Z(
        mux_b[6]) );
  LVT_AO22HSV2 U28 ( .A1(mux_bq[7]), .A2(n11), .B1(b_out[7]), .B2(n18), .Z(
        mux_b[7]) );
  LVT_AO22HSV4 U29 ( .A1(ti_7[2]), .A2(ctro), .B1(t_i_2_out[2]), .B2(n20), .Z(
        to_7[2]) );
  LVT_AO22HSV4 U30 ( .A1(ti_7[3]), .A2(ctro), .B1(t_i_2_out[3]), .B2(n20), .Z(
        to_7[3]) );
  LVT_AO22HSV4 U31 ( .A1(ti_7[4]), .A2(ctro), .B1(t_i_2_out[4]), .B2(n20), .Z(
        to_7[4]) );
  LVT_AO22HSV4 U32 ( .A1(ti_7[6]), .A2(ctro), .B1(t_i_2_out[6]), .B2(n20), .Z(
        to_7[6]) );
  LVT_MOAI22HSV4 U33 ( .A1(l_ctr), .A2(n19), .B1(ti_1), .B2(l_ctr), .ZN(to_1)
         );
  LVT_INHSV2 U34 ( .I(rstn), .ZN(n15) );
endmodule


module regist_8bit_95 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_94 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_93 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_63 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_62 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_63 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV4 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV4 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV4 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_62 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
endmodule


module regist_1bit_61 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_92 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_60 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_61 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module cell_3_799 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_111 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_110 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_109 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_108 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_107 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV2 U1 ( .A1(n5), .A2(n2), .A3(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_106 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XNOR2HSV1 U1 ( .A1(n1), .A2(n7), .ZN(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV1 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n1) );
endmodule


module cell_4_105 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n9) );
  LVT_INAND2HSV0 U1 ( .A1(n9), .B1(n8), .ZN(n5) );
  LVT_CLKNHSV2 U2 ( .I(n8), .ZN(n1) );
  LVT_CLKNAND2HSV2 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n1), .A2(n9), .ZN(n6) );
  LVT_NAND2HSV2 U6 ( .A1(n5), .A2(n6), .ZN(n10) );
  LVT_XNOR2HSV4 U7 ( .A1(n10), .A2(n7), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U8 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_1_15 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_3_799 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_111 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(
        t_i_1_out[1]) );
  cell_4_110 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_109 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(
        t_i_1_out[3]) );
  cell_4_108 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(t_i_1_out[4])
         );
  cell_4_107 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(
        t_i_1_out[5]) );
  cell_4_106 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_105 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_111 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_798 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_797 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_796 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_795 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_794 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_793 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_792 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n9) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_OAI21HSV2 U2 ( .A1(n10), .A2(n8), .B(n2), .ZN(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(n10), .A2(n8), .ZN(n2) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U6 ( .A1(t_i_1_in), .A2(n9), .ZN(n6) );
  LVT_CLKNHSV2 U7 ( .I(t_i_1_in), .ZN(n4) );
  LVT_NAND2HSV2 U8 ( .A1(n6), .A2(n7), .ZN(n8) );
  LVT_INHSV2 U9 ( .I(n9), .ZN(n5) );
endmodule


module row_other_111 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_111 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_798 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_797 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_796 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_795 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_794 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_793 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_792 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_110 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_791 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_790 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_789 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_788 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_787 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_786 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(g_in), .A2(t_m_1_in), .ZN(n6) );
endmodule


module cell_3_785 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U2 ( .A1(n8), .A2(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV2 U4 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV2 U5 ( .A1(n5), .A2(n6), .ZN(n7) );
  LVT_INHSV2 U6 ( .I(n8), .ZN(n2) );
  LVT_INHSV2 U7 ( .I(t_i_1_in), .ZN(n4) );
  LVT_XNOR2HSV4 U8 ( .A1(n9), .A2(n7), .ZN(t_i_out) );
endmodule


module row_other_110 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_110 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_791 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_790 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_789 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_788 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_787 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_786 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_785 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_109 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_784 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_783 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_782 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_781 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_780 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_XNOR2HSV1 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_779 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV1 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module cell_3_778 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XNOR2HSV1 U1 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U4 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U6 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV2 U7 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV1 U8 ( .A1(n9), .A2(n7), .ZN(n5) );
endmodule


module row_other_109 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_109 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_784 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_783 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_782 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_781 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_780 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_779 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_778 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_108 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_777 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_776 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_775 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_774 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_773 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_772 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_771 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U2 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U5 ( .I(n7), .ZN(n4) );
  LVT_INHSV2SR U6 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV0P5 U7 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_108 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_108 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_777 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_776 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_775 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_774 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_773 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_772 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_771 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_107 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_770 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_769 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_768 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_767 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_766 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV1 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_765 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_764 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .Z(n3) );
  LVT_XOR2HSV4 U3 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n3), .A2(t_i_1_in), .ZN(n4) );
endmodule


module row_other_107 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_107 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_770 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_769 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_768 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_767 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_766 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_765 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_764 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_106 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n3), .A2(n4), .Z(t_i_out) );
endmodule


module cell_3_763 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_XNOR2HSV1 U1 ( .A1(t_i_1_in), .A2(n3), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U3 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_CLKAND2HSV2 U4 ( .A1(b_in), .A2(a_in), .Z(n3) );
endmodule


module cell_3_762 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_761 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_760 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_759 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_758 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_757 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV4SR U2 ( .I(n9), .ZN(n2) );
  LVT_CLKNHSV4 U4 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV4 U5 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U7 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_106 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_106 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_763 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_762 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_761 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_760 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_759 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_758 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_757 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_105 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n3), .A2(n4), .Z(t_i_out) );
endmodule


module cell_3_756 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_755 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U2 ( .A1(t_i_1_in), .A2(n4), .ZN(n5) );
  LVT_INHSV2 U4 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV1 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XOR2HSV0 U6 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_3_754 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_INHSV2SR U4 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_XOR2HSV2 U6 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
endmodule


module cell_3_753 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n12) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n14) );
  LVT_NAND2HSV1 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNHSV0 U4 ( .I(n14), .ZN(n8) );
  LVT_NAND2HSV2 U5 ( .A1(n12), .A2(n5), .ZN(n6) );
  LVT_CLKNAND2HSV1 U6 ( .A1(n6), .A2(n7), .ZN(n13) );
  LVT_INHSV2 U7 ( .I(n12), .ZN(n4) );
  LVT_INHSV2 U8 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV0 U9 ( .A1(n9), .A2(n14), .ZN(n10) );
  LVT_NAND2HSV0P5 U10 ( .A1(n8), .A2(n13), .ZN(n11) );
  LVT_NAND2HSV1 U11 ( .A1(n10), .A2(n11), .ZN(t_i_out) );
  LVT_CLKNHSV1 U12 ( .I(n13), .ZN(n9) );
endmodule


module cell_3_752 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_751 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_XNOR2HSV1 U1 ( .A1(t_i_1_in), .A2(n3), .ZN(n4) );
  LVT_CLKAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .Z(n3) );
  LVT_NAND2HSV1 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n5), .A2(n4), .Z(t_i_out) );
endmodule


module cell_3_750 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module row_other_105 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_105 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_756 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_755 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_754 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_753 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_752 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_751 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_750 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_15 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_15 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(
        t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), 
        .t_i_1_out(t0), .t_i_2_out(t_i_2_out[6]) );
  row_other_111 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_110 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_109 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_108 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_107 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_106 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_105 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_91 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_90 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_7bit_60 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module PE_15 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, 
        t_i_2_in, a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro
 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  LVT_AO22HSV0 U15 ( .A1(mux_bq[3]), .A2(n15), .B1(b_out[3]), .B2(n12), .Z(
        mux_b[3]) );
  LVT_AO22HSV0 U16 ( .A1(mux_bq[2]), .A2(n15), .B1(b_out[2]), .B2(n12), .Z(
        mux_b[2]) );
  LVT_AO22HSV0 U17 ( .A1(mux_bq[1]), .A2(n15), .B1(b_out[1]), .B2(n12), .Z(
        mux_b[1]) );
  regist_8bit_95 u0 ( .clk(clk), .rstn(n18), .in(a_in), .out(l_a) );
  regist_8bit_94 u1 ( .clk(clk), .rstn(n18), .in(b_in), .out(b_out) );
  regist_8bit_93 u2 ( .clk(clk), .rstn(n18), .in(g_in), .out(l_g) );
  regist_1bit_63 u3 ( .clk(clk), .rstn(n18), .in(ctr), .out(l_ctr) );
  regist_1bit_62 u4 ( .clk(clk), .rstn(n18), .in(n15), .out(ctro) );
  regist_7bit_63 u5 ( .clk(clk), .rstn(n18), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_7bit_62 u6 ( .clk(clk), .rstn(n18), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_61 u7 ( .clk(clk), .rstn(n18), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_8bit_92 u9 ( .clk(clk), .rstn(n18), .in(mux_b), .out(mux_bq) );
  regist_1bit_60 u10 ( .clk(clk), .rstn(n18), .in(n14), .out(ti_1) );
  regist_7bit_61 u11 ( .clk(clk), .rstn(n18), .in(to_7), .out(ti_7) );
  PE_core_15 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out(t_i_2_out), .t_i_1_out_0(t_i_1_out_0)
         );
  regist_8bit_91 u12 ( .clk(clk), .rstn(n18), .in(ao), .out(a_out) );
  regist_8bit_90 u13 ( .clk(clk), .rstn(n18), .in(go), .out(g_out) );
  regist_7bit_60 u14 ( .clk(clk), .rstn(n18), .in(to), .out(t_i_1_out) );
  LVT_NOR2HSV1 U2 ( .A1(n23), .A2(n22), .ZN(c_t_i_1_in_0) );
  LVT_AOI21HSV2 U3 ( .A1(n21), .A2(n20), .B(n22), .ZN(\c_t_i_1_in[0] ) );
  LVT_INHSV2 U4 ( .I(ctro), .ZN(n24) );
  LVT_NAND2HSV2 U5 ( .A1(ti_7[1]), .A2(ctro), .ZN(n16) );
  LVT_NOR3HSV2 U6 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), 
        .ZN(n21) );
  LVT_CLKNAND2HSV4 U7 ( .A1(n6), .A2(n7), .ZN(to_7[3]) );
  LVT_CLKNAND2HSV8 U8 ( .A1(n17), .A2(n16), .ZN(to_7[1]) );
  LVT_NAND2HSV2 U9 ( .A1(ti_7[3]), .A2(ctro), .ZN(n6) );
  LVT_CLKNAND2HSV3 U10 ( .A1(t_i_2_out[3]), .A2(n24), .ZN(n7) );
  LVT_NAND2HSV2 U11 ( .A1(ti_7[2]), .A2(ctro), .ZN(n8) );
  LVT_CLKNAND2HSV2 U12 ( .A1(t_i_2_out[2]), .A2(n24), .ZN(n9) );
  LVT_NAND2HSV4 U13 ( .A1(n8), .A2(n9), .ZN(to_7[2]) );
  LVT_CLKNAND2HSV3 U14 ( .A1(ti_7[5]), .A2(ctro), .ZN(n10) );
  LVT_CLKNAND2HSV3 U18 ( .A1(t_i_2_out[5]), .A2(n24), .ZN(n11) );
  LVT_NAND2HSV4 U19 ( .A1(n10), .A2(n11), .ZN(to_7[5]) );
  LVT_NAND2HSV4 U20 ( .A1(t_i_2_out[1]), .A2(n24), .ZN(n17) );
  LVT_INHSV4SR U21 ( .I(l_t_i_1_in_0), .ZN(n23) );
  LVT_INHSV6 U22 ( .I(n19), .ZN(n18) );
  LVT_BUFHSV2RT U23 ( .I(n22), .Z(n12) );
  LVT_INHSV0SR U24 ( .I(l_ctr), .ZN(n22) );
  LVT_INHSV0SR U25 ( .I(to_1), .ZN(n13) );
  LVT_INHSV2 U26 ( .I(n13), .ZN(n14) );
  LVT_NOR4HSV12 U27 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(
        l_t_i_1_in[4]), .A4(l_t_i_1_in[3]), .ZN(n20) );
  LVT_INHSV2 U28 ( .I(n22), .ZN(n15) );
  LVT_AO22HSV2 U29 ( .A1(mux_bq[4]), .A2(n15), .B1(b_out[4]), .B2(n12), .Z(
        mux_b[4]) );
  LVT_AO22HSV2 U30 ( .A1(mux_bq[0]), .A2(n15), .B1(b_out[0]), .B2(n12), .Z(
        mux_b[0]) );
  LVT_AO22HSV2 U31 ( .A1(mux_bq[6]), .A2(n15), .B1(b_out[6]), .B2(n12), .Z(
        mux_b[6]) );
  LVT_AO22HSV2 U32 ( .A1(mux_bq[7]), .A2(n15), .B1(b_out[7]), .B2(n12), .Z(
        mux_b[7]) );
  LVT_AO22HSV2 U33 ( .A1(mux_bq[5]), .A2(n15), .B1(b_out[5]), .B2(n12), .Z(
        mux_b[5]) );
  LVT_AO22HSV4 U34 ( .A1(ti_7[0]), .A2(ctro), .B1(t_i_2_out[0]), .B2(n24), .Z(
        to_7[0]) );
  LVT_AO22HSV4 U35 ( .A1(ti_7[4]), .A2(ctro), .B1(t_i_2_out[4]), .B2(n24), .Z(
        to_7[4]) );
  LVT_AO22HSV4 U36 ( .A1(ti_7[6]), .A2(ctro), .B1(t_i_2_out[6]), .B2(n24), .Z(
        to_7[6]) );
  LVT_MOAI22HSV4 U37 ( .A1(l_ctr), .A2(n23), .B1(l_ctr), .B2(ti_1), .ZN(to_1)
         );
  LVT_INHSV2 U38 ( .I(rstn), .ZN(n19) );
endmodule


module regist_8bit_89 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_88 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_87 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_59 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_58 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_59 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV4 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV4 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV4 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_58 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
endmodule


module regist_1bit_57 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_86 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_56 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_57 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module cell_3_749 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_104 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_103 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_102 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U3 ( .A1(n6), .A2(n5), .Z(n7) );
endmodule


module cell_4_101 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_100 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_XOR2HSV2 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_99 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV2 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_98 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n13) );
  LVT_INAND2HSV0 U1 ( .A1(n13), .B1(n12), .ZN(n10) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n12) );
  LVT_NAND2HSV1 U3 ( .A1(n11), .A2(n14), .ZN(n6) );
  LVT_XNOR2HSV1 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n11) );
  LVT_NAND2HSV4 U6 ( .A1(n1), .A2(n5), .ZN(n7) );
  LVT_CLKNHSV0P5 U7 ( .I(n12), .ZN(n8) );
  LVT_CLKNAND2HSV2 U8 ( .A1(n8), .A2(n13), .ZN(n9) );
  LVT_INHSV2 U9 ( .I(n14), .ZN(n1) );
  LVT_CLKNAND2HSV3 U10 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV3SR U11 ( .I(n11), .ZN(n5) );
  LVT_NAND2HSV2 U12 ( .A1(n9), .A2(n10), .ZN(n14) );
endmodule


module row_1_14 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_3_749 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_104 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(
        t_i_1_out[1]) );
  cell_4_103 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_102 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(
        t_i_1_out[3]) );
  cell_4_101 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(
        t_i_1_out[4]) );
  cell_4_100 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(
        t_i_1_out[5]) );
  cell_4_99 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_98 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_104 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_748 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_747 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_746 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_745 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_744 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_743 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV2 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_742 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U4 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV3 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV2 U6 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV0 U7 ( .A1(n7), .A2(n9), .ZN(n5) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_104 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_104 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_748 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_747 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_746 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_745 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_744 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_743 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_742 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_103 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_741 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_740 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_739 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_738 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_737 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_736 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_735 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4;

  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U2 ( .A1(t_i_1_in), .A2(n2), .Z(n3) );
  LVT_CLKAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .Z(n2) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(n3), .ZN(t_i_out) );
endmodule


module row_other_103 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_103 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_741 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_740 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_739 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_738 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_737 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_736 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_735 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_102 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_734 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_733 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_732 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_731 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_730 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_729 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_728 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV3SR U1 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV3 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV0P5 U4 ( .A1(n7), .A2(n9), .ZN(n5) );
  LVT_INHSV3 U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV4 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_102 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_102 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_734 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_733 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_732 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_731 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_730 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_729 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_728 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2SR U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_101 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n3), .A2(n4), .Z(t_i_out) );
endmodule


module cell_3_727 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_726 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_725 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_724 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_723 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_722 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV2 U4 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U5 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV0P5 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2SR U7 ( .I(n9), .ZN(n2) );
  LVT_INHSV2 U8 ( .I(n7), .ZN(n4) );
endmodule


module cell_3_721 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  LVT_CLKNAND2HSV3 U1 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_CLKNHSV0P5 U2 ( .I(n13), .ZN(n5) );
  LVT_NAND2HSV2 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n14) );
  LVT_INHSV2 U4 ( .I(n14), .ZN(n4) );
  LVT_NAND2HSV2 U5 ( .A1(n10), .A2(n11), .ZN(n13) );
  LVT_NAND2HSV2 U6 ( .A1(n12), .A2(n9), .ZN(n10) );
  LVT_CLKNAND2HSV1 U7 ( .A1(n14), .A2(n5), .ZN(n6) );
  LVT_INHSV2 U8 ( .I(t_i_1_in), .ZN(n9) );
  LVT_NAND2HSV4 U9 ( .A1(n4), .A2(n13), .ZN(n7) );
  LVT_NAND2HSV2 U10 ( .A1(n8), .A2(t_i_1_in), .ZN(n11) );
  LVT_INHSV2 U11 ( .I(n12), .ZN(n8) );
  LVT_NAND2HSV0 U12 ( .A1(b_in), .A2(a_in), .ZN(n12) );
endmodule


module row_other_101 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_101 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_727 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_726 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_725 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_724 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_723 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_722 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_721 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_100 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_720 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_719 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_718 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_717 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_716 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_715 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_714 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV2 U2 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV2 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2 U5 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_100 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_100 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_720 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_719 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_718 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_717 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_716 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_715 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_714 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_99 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_713 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_712 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_711 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_710 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_709 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_708 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_707 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV3SR U2 ( .I(n9), .ZN(n2) );
  LVT_INHSV3 U4 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n7), .A2(n9), .ZN(n5) );
  LVT_NAND2HSV4 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_99 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_99 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_713 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_712 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_711 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_710 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_709 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_708 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_707 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_98 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_706 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_INAND2HSV0 U1 ( .A1(n8), .B1(n9), .ZN(n5) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XOR2HSV0 U4 ( .A1(t_i_1_in), .A2(n7), .Z(n8) );
  LVT_CLKNAND2HSV0 U5 ( .A1(n4), .A2(n8), .ZN(n6) );
  LVT_NAND2HSV0 U6 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV0P5SR U7 ( .I(n9), .ZN(n4) );
endmodule


module cell_3_705 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_704 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_703 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_702 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKXOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_701 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_700 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module row_other_98 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_98 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_706 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_705 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_704 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_703 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_702 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_701 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_700 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_14 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_14 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(
        t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), 
        .t_i_1_out(t0), .t_i_2_out(t_i_2_out[6]) );
  row_other_104 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_103 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_102 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_101 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_100 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_99 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_98 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_85 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_84 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_7bit_56 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
endmodule


module PE_14 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, 
        t_i_2_in, a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro
 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1, n3,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  regist_8bit_89 u0 ( .clk(clk), .rstn(n12), .in(a_in), .out(l_a) );
  regist_8bit_88 u1 ( .clk(clk), .rstn(n12), .in(b_in), .out(b_out) );
  regist_8bit_87 u2 ( .clk(clk), .rstn(n12), .in(g_in), .out(l_g) );
  regist_1bit_59 u3 ( .clk(clk), .rstn(n12), .in(ctr), .out(l_ctr) );
  regist_1bit_58 u4 ( .clk(clk), .rstn(n12), .in(n11), .out(ctro) );
  regist_7bit_59 u5 ( .clk(clk), .rstn(n12), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_7bit_58 u6 ( .clk(clk), .rstn(n12), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_57 u7 ( .clk(clk), .rstn(n12), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_8bit_86 u9 ( .clk(clk), .rstn(n12), .in(mux_b), .out(mux_bq) );
  regist_1bit_56 u10 ( .clk(clk), .rstn(n12), .in(n9), .out(ti_1) );
  regist_7bit_57 u11 ( .clk(clk), .rstn(n12), .in(to_7), .out(ti_7) );
  PE_core_14 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out(t_i_2_out), .t_i_1_out_0(t_i_1_out_0)
         );
  regist_8bit_85 u12 ( .clk(clk), .rstn(n12), .in(ao), .out(a_out) );
  regist_8bit_84 u13 ( .clk(clk), .rstn(n12), .in(go), .out(g_out) );
  regist_7bit_56 u14 ( .clk(clk), .rstn(n12), .in(to), .out(t_i_1_out) );
  LVT_CLKNAND2HSV8 U2 ( .A1(n7), .A2(n8), .ZN(to_7[2]) );
  LVT_INHSV2P5 U3 ( .I(l_ctr), .ZN(n10) );
  LVT_INHSV2 U4 ( .I(ctro), .ZN(n17) );
  LVT_NAND2HSV4 U5 ( .A1(t_i_2_out[2]), .A2(n17), .ZN(n8) );
  LVT_AO22HSV1 U6 ( .A1(mux_bq[5]), .A2(n11), .B1(b_out[5]), .B2(n10), .Z(
        mux_b[5]) );
  LVT_AO22HSV1 U7 ( .A1(mux_bq[7]), .A2(n11), .B1(b_out[7]), .B2(n10), .Z(
        mux_b[7]) );
  LVT_AO22HSV1 U8 ( .A1(mux_bq[6]), .A2(n11), .B1(b_out[6]), .B2(n10), .Z(
        mux_b[6]) );
  LVT_AO22HSV1 U9 ( .A1(mux_bq[3]), .A2(n11), .B1(b_out[3]), .B2(n10), .Z(
        mux_b[3]) );
  LVT_AO22HSV1 U10 ( .A1(mux_bq[2]), .A2(n11), .B1(b_out[2]), .B2(n10), .Z(
        mux_b[2]) );
  LVT_AO22HSV1 U11 ( .A1(mux_bq[0]), .A2(n11), .B1(b_out[0]), .B2(n10), .Z(
        mux_b[0]) );
  LVT_NOR3HSV2 U12 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), .ZN(n15) );
  LVT_INHSV4 U13 ( .I(l_t_i_1_in_0), .ZN(n16) );
  LVT_NAND2HSV2 U14 ( .A1(ti_7[6]), .A2(ctro), .ZN(n3) );
  LVT_CLKNAND2HSV4 U15 ( .A1(t_i_2_out[6]), .A2(n17), .ZN(n6) );
  LVT_NAND2HSV4 U16 ( .A1(n3), .A2(n6), .ZN(to_7[6]) );
  LVT_NAND2HSV2 U17 ( .A1(ti_7[2]), .A2(ctro), .ZN(n7) );
  LVT_INHSV6 U18 ( .I(n13), .ZN(n12) );
  LVT_IOA22HSV0 U19 ( .B1(l_ctr), .B2(n16), .A1(ti_1), .A2(l_ctr), .ZN(n9) );
  LVT_MOAI22HSV4 U20 ( .A1(n16), .A2(l_ctr), .B1(l_ctr), .B2(ti_1), .ZN(to_1)
         );
  LVT_NOR2HSV0 U21 ( .A1(n16), .A2(n10), .ZN(c_t_i_1_in_0) );
  LVT_NOR4HSV12 U22 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(
        l_t_i_1_in[4]), .A4(l_t_i_1_in[3]), .ZN(n14) );
  LVT_INHSV2 U23 ( .I(n10), .ZN(n11) );
  LVT_AOI21HSV1 U24 ( .A1(n15), .A2(n14), .B(n10), .ZN(\c_t_i_1_in[0] ) );
  LVT_AO22HSV2 U25 ( .A1(mux_bq[1]), .A2(n11), .B1(b_out[1]), .B2(n10), .Z(
        mux_b[1]) );
  LVT_AO22HSV2 U26 ( .A1(mux_bq[4]), .A2(n11), .B1(b_out[4]), .B2(n10), .Z(
        mux_b[4]) );
  LVT_AO22HSV4 U27 ( .A1(ti_7[0]), .A2(ctro), .B1(t_i_2_out[0]), .B2(n17), .Z(
        to_7[0]) );
  LVT_AO22HSV4 U28 ( .A1(ti_7[1]), .A2(ctro), .B1(t_i_2_out[1]), .B2(n17), .Z(
        to_7[1]) );
  LVT_AO22HSV4 U29 ( .A1(ti_7[3]), .A2(ctro), .B1(t_i_2_out[3]), .B2(n17), .Z(
        to_7[3]) );
  LVT_AO22HSV4 U30 ( .A1(ti_7[4]), .A2(ctro), .B1(t_i_2_out[4]), .B2(n17), .Z(
        to_7[4]) );
  LVT_AO22HSV4 U31 ( .A1(ti_7[5]), .A2(ctro), .B1(t_i_2_out[5]), .B2(n17), .Z(
        to_7[5]) );
  LVT_INHSV2 U32 ( .I(rstn), .ZN(n13) );
endmodule


module regist_8bit_83 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_82 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_81 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_55 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_54 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV1 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_55 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV4 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV4 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV4 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV4 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV4 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_54 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
endmodule


module regist_1bit_53 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_80 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_52 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_53 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module cell_3_699 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_97 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV2 U5 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_96 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_95 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_94 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n5, n6, n7, n8, n9, n10, n11;

  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n11) );
  LVT_CLKNHSV2 U1 ( .I(n9), .ZN(n5) );
  LVT_XNOR2HSV1 U2 ( .A1(n11), .A2(n8), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV0 U4 ( .A1(n10), .A2(n9), .ZN(n6) );
  LVT_NAND2HSV0P5 U6 ( .A1(n2), .A2(n5), .ZN(n7) );
  LVT_NAND2HSV2 U7 ( .A1(n6), .A2(n7), .ZN(n8) );
  LVT_CLKNHSV2 U8 ( .I(n10), .ZN(n2) );
  LVT_NAND2HSV2 U9 ( .A1(b_in), .A2(a_in), .ZN(n10) );
endmodule


module cell_4_93 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n5, n6, n7;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n7) );
  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(n2) );
  LVT_XOR2HSV2 U2 ( .A1(n7), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_92 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n2, n4;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR3HSV2 U1 ( .A1(n1), .A2(n2), .A3(n4), .ZN(t_i_out) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_XNOR2HSV1 U3 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n1) );
endmodule


module cell_4_91 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n5, n6, n7;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n7) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n7), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U3 ( .A1(n5), .A2(n6), .ZN(n2) );
endmodule


module row_1_13 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_3_699 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_97 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(
        t_i_1_out[1]) );
  cell_4_96 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_95 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(
        t_i_1_out[3]) );
  cell_4_94 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(
        t_i_1_out[4]) );
  cell_4_93 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(
        t_i_1_out[5]) );
  cell_4_92 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_91 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_97 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_698 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_697 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_CLKAND2HSV2 U1 ( .A1(b_in), .A2(a_in), .Z(n3) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U3 ( .A1(n3), .A2(t_i_1_in), .ZN(n4) );
  LVT_XOR2HSV2 U4 ( .A1(n5), .A2(n4), .Z(t_i_out) );
endmodule


module cell_3_696 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_695 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_694 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_693 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV2 U5 ( .I(n8), .ZN(n4) );
  LVT_INHSV2 U6 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV2 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_XOR2HSV2 U8 ( .A1(n10), .A2(n9), .Z(t_i_out) );
endmodule


module cell_3_692 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n6), .Z(n7) );
  LVT_CLKAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .Z(n6) );
  LVT_INHSV2 U3 ( .I(n7), .ZN(n3) );
  LVT_CLKNAND2HSV0 U4 ( .A1(n8), .A2(n7), .ZN(n4) );
  LVT_CLKNAND2HSV3 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_NAND2HSV4 U6 ( .A1(n2), .A2(n3), .ZN(n5) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n4), .A2(n5), .ZN(t_i_out) );
  LVT_INHSV3SR U8 ( .I(n8), .ZN(n2) );
endmodule


module row_other_97 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_97 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_698 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_697 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_696 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_695 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_694 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_693 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_692 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_96 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_691 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_690 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_689 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_688 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module cell_3_687 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_686 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module cell_3_685 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_96 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_96 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_691 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_690 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_689 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_688 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_687 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_686 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_685 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_95 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_684 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_683 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_682 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_681 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_680 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_679 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_678 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNHSV2 U2 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV2 U4 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV1 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV3 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_95 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_95 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_684 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_683 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_682 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_681 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_680 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_679 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_678 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_94 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_677 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_676 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_675 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_674 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_673 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_672 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_671 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n2), .A2(n6), .ZN(n5) );
  LVT_NAND2HSV3 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNHSV2 U4 ( .I(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U6 ( .A1(t_i_1_in), .A2(n8), .ZN(n4) );
  LVT_INHSV2 U7 ( .I(n8), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(n9), .A2(n7), .ZN(t_i_out) );
endmodule


module row_other_94 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_94 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_677 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_676 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_675 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_674 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_673 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_672 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_671 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_93 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n3), .A2(n4), .Z(t_i_out) );
endmodule


module cell_3_670 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_669 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_668 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_667 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_666 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_665 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_XNOR2HSV1 U1 ( .A1(t_i_1_in), .A2(n3), .ZN(n4) );
  LVT_CLKAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .Z(n3) );
  LVT_CLKXOR2HSV4 U3 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_664 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U5 ( .I(n9), .ZN(n2) );
  LVT_INHSV2 U6 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV0P5 U7 ( .A1(n7), .A2(n9), .ZN(n5) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_93 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_93 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_670 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_669 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_668 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_667 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_666 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_665 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_664 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_92 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_663 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_662 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_661 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_660 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_659 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_658 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U4 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_INHSV0SR U6 ( .I(n8), .ZN(n4) );
endmodule


module cell_3_657 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2SR U5 ( .I(n9), .ZN(n2) );
  LVT_CLKNHSV5 U6 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV4 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_92 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_92 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_663 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_662 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_661 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_660 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_659 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_658 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_657 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_91 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n3), .A2(n4), .Z(t_i_out) );
endmodule


module cell_3_656 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_655 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_654 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_653 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_652 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_651 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_650 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module row_other_91 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_91 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_656 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_655 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_654 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_653 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_652 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_651 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_650 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_13 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_13 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(
        t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), 
        .t_i_1_out(t0), .t_i_2_out(t_i_2_out[6]) );
  row_other_97 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_96 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_95 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_94 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_93 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_92 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_91 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_79 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_78 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_7bit_52 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
endmodule


module PE_13 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, 
        t_i_2_in, a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro
 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  LVT_NOR3HSV0 U24 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), .ZN(n16) );
  regist_8bit_83 u0 ( .clk(clk), .rstn(n13), .in(a_in), .out(l_a) );
  regist_8bit_82 u1 ( .clk(clk), .rstn(n13), .in(b_in), .out(b_out) );
  regist_8bit_81 u2 ( .clk(clk), .rstn(n13), .in(g_in), .out(l_g) );
  regist_1bit_55 u3 ( .clk(clk), .rstn(n13), .in(ctr), .out(l_ctr) );
  regist_1bit_54 u4 ( .clk(clk), .rstn(n13), .in(n8), .out(ctro) );
  regist_7bit_55 u5 ( .clk(clk), .rstn(n13), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_7bit_54 u6 ( .clk(clk), .rstn(n13), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_53 u7 ( .clk(clk), .rstn(n13), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_8bit_80 u9 ( .clk(clk), .rstn(n13), .in(mux_b), .out(mux_bq) );
  regist_1bit_52 u10 ( .clk(clk), .rstn(n13), .in(to_1), .out(ti_1) );
  regist_7bit_53 u11 ( .clk(clk), .rstn(n13), .in(to_7), .out(ti_7) );
  PE_core_13 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out(t_i_2_out), .t_i_1_out_0(t_i_1_out_0)
         );
  regist_8bit_79 u12 ( .clk(clk), .rstn(n13), .in(ao), .out(a_out) );
  regist_8bit_78 u13 ( .clk(clk), .rstn(n13), .in(go), .out(g_out) );
  regist_7bit_52 u14 ( .clk(clk), .rstn(n13), .in(to), .out(t_i_1_out) );
  LVT_NOR2HSV1 U2 ( .A1(n18), .A2(n17), .ZN(c_t_i_1_in_0) );
  LVT_INHSV2 U3 ( .I(l_ctr), .ZN(n17) );
  LVT_INHSV4SR U4 ( .I(l_t_i_1_in_0), .ZN(n18) );
  LVT_NAND2HSV2 U5 ( .A1(ti_7[6]), .A2(ctro), .ZN(n11) );
  LVT_NAND2HSV4 U6 ( .A1(t_i_2_out[6]), .A2(n19), .ZN(n12) );
  LVT_AO22HSV1 U7 ( .A1(mux_bq[2]), .A2(n8), .B1(b_out[2]), .B2(n17), .Z(
        mux_b[2]) );
  LVT_AO22HSV1 U8 ( .A1(mux_bq[6]), .A2(n8), .B1(b_out[6]), .B2(n17), .Z(
        mux_b[6]) );
  LVT_AO22HSV1 U9 ( .A1(mux_bq[7]), .A2(n8), .B1(b_out[7]), .B2(n17), .Z(
        mux_b[7]) );
  LVT_AO22HSV1 U10 ( .A1(mux_bq[0]), .A2(n8), .B1(b_out[0]), .B2(n17), .Z(
        mux_b[0]) );
  LVT_AO22HSV1 U11 ( .A1(mux_bq[1]), .A2(n8), .B1(b_out[1]), .B2(n17), .Z(
        mux_b[1]) );
  LVT_NAND2HSV2 U12 ( .A1(ti_7[4]), .A2(ctro), .ZN(n9) );
  LVT_NAND2HSV4 U13 ( .A1(t_i_2_out[4]), .A2(n19), .ZN(n10) );
  LVT_CLKNAND2HSV1 U14 ( .A1(ti_7[2]), .A2(ctro), .ZN(n6) );
  LVT_NAND2HSV4 U15 ( .A1(t_i_2_out[2]), .A2(n19), .ZN(n7) );
  LVT_NAND2HSV8 U16 ( .A1(n6), .A2(n7), .ZN(to_7[2]) );
  LVT_INHSV2 U17 ( .I(ctro), .ZN(n19) );
  LVT_INHSV6 U18 ( .I(n14), .ZN(n13) );
  LVT_NOR4HSV12 U19 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(
        l_t_i_1_in[4]), .A4(l_t_i_1_in[3]), .ZN(n15) );
  LVT_BUFHSV2RT U20 ( .I(l_ctr), .Z(n8) );
  LVT_CLKNAND2HSV8 U21 ( .A1(n10), .A2(n9), .ZN(to_7[4]) );
  LVT_CLKNAND2HSV8 U22 ( .A1(n12), .A2(n11), .ZN(to_7[6]) );
  LVT_AOI21HSV2 U23 ( .A1(n16), .A2(n15), .B(n17), .ZN(\c_t_i_1_in[0] ) );
  LVT_AO22HSV2 U25 ( .A1(mux_bq[3]), .A2(n8), .B1(b_out[3]), .B2(n17), .Z(
        mux_b[3]) );
  LVT_AO22HSV2 U26 ( .A1(mux_bq[4]), .A2(n8), .B1(b_out[4]), .B2(n17), .Z(
        mux_b[4]) );
  LVT_AO22HSV2 U27 ( .A1(mux_bq[5]), .A2(n8), .B1(b_out[5]), .B2(n17), .Z(
        mux_b[5]) );
  LVT_AO22HSV4 U28 ( .A1(ti_7[0]), .A2(ctro), .B1(t_i_2_out[0]), .B2(n19), .Z(
        to_7[0]) );
  LVT_AO22HSV4 U29 ( .A1(ti_7[1]), .A2(ctro), .B1(t_i_2_out[1]), .B2(n19), .Z(
        to_7[1]) );
  LVT_AO22HSV4 U30 ( .A1(ti_7[3]), .A2(ctro), .B1(t_i_2_out[3]), .B2(n19), .Z(
        to_7[3]) );
  LVT_AO22HSV4 U31 ( .A1(ti_7[5]), .A2(ctro), .B1(t_i_2_out[5]), .B2(n19), .Z(
        to_7[5]) );
  LVT_MOAI22HSV4 U32 ( .A1(n18), .A2(l_ctr), .B1(ti_1), .B2(l_ctr), .ZN(to_1)
         );
  LVT_INHSV2 U33 ( .I(rstn), .ZN(n14) );
endmodule


module regist_8bit_77 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_76 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_75 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_51 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_50 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_51 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_50 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
endmodule


module regist_1bit_49 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_74 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_48 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_49 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module cell_3_649 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_90 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U3 ( .A1(t_i_1_in), .A2(t_i_2_in), .Z(n8) );
  LVT_XOR2HSV0 U5 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_89 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_88 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_XOR3HSV1 U2 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
endmodule


module cell_4_87 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n2), .A3(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_86 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_XOR3HSV1 U2 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
endmodule


module cell_4_85 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U3 ( .A1(n6), .A2(n5), .Z(n7) );
endmodule


module cell_4_84 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n6), .A2(n7), .Z(n8) );
  LVT_OAI21HSV2 U3 ( .A1(n5), .A2(n8), .B(n1), .ZN(t_i_out) );
  LVT_NAND2HSV2 U5 ( .A1(n5), .A2(n8), .ZN(n1) );
  LVT_XNOR2HSV1 U6 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n5) );
endmodule


module row_1_12 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_3_649 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_90 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(
        t_i_1_out[1]) );
  cell_4_89 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_88 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(t_i_1_out[3])
         );
  cell_4_87 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(
        t_i_1_out[4]) );
  cell_4_86 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(t_i_1_out[5])
         );
  cell_4_85 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_84 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U3 ( .I(n2), .ZN(n3) );
  LVT_CLKNHSV0P5 U4 ( .I(n3), .ZN(n4) );
endmodule


module cell_2_90 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_648 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_647 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_646 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_645 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_644 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_643 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV2 U3 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U4 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV2 U5 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV1 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_642 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;

  LVT_NAND2HSV2 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV2 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n13) );
  LVT_NAND2HSV2 U4 ( .A1(n9), .A2(n10), .ZN(n11) );
  LVT_INHSV2SR U5 ( .I(n13), .ZN(n2) );
  LVT_CLKNAND2HSV0 U6 ( .A1(n13), .A2(n11), .ZN(n5) );
  LVT_INHSV2SR U7 ( .I(n11), .ZN(n4) );
  LVT_CLKNHSV2 U8 ( .I(t_i_1_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U9 ( .A1(n12), .A2(t_i_1_in), .ZN(n9) );
  LVT_CLKNAND2HSV1 U10 ( .A1(n7), .A2(n8), .ZN(n10) );
  LVT_INHSV2 U11 ( .I(n12), .ZN(n7) );
  LVT_NAND2HSV0 U12 ( .A1(b_in), .A2(a_in), .ZN(n12) );
endmodule


module row_other_90 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_90 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_648 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_647 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_646 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_645 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_644 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_643 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_642 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_89 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_641 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_640 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_639 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_638 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_637 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_636 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_635 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U1 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2 U2 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U4 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNAND2HSV3 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV2 U6 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV4 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U8 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
endmodule


module row_other_89 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_89 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_641 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_640 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_639 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_638 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_637 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_636 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_635 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_88 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_634 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_633 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_632 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_631 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_630 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_629 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_628 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV2 U1 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2SR U4 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV2 U5 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV2 U7 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV2 U8 ( .A1(n9), .A2(n7), .ZN(n5) );
endmodule


module row_other_88 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_88 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_634 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_633 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_632 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_631 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_630 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_629 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_628 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_87 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_627 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_626 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_625 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_624 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_623 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_622 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_621 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module row_other_87 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_87 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_627 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_626 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_625 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_624 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_623 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_622 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_621 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_86 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n3), .A2(n4), .Z(t_i_out) );
endmodule


module cell_3_620 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_619 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_618 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_617 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_616 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_615 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_614 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV2 U2 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNHSV4 U4 ( .I(n7), .ZN(n4) );
  LVT_INHSV2 U5 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV0P5 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV4 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U8 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
endmodule


module row_other_86 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_86 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_620 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_619 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_618 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_617 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_616 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_615 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_614 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_85 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_613 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_612 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_611 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_610 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_609 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_608 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_607 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV4 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNHSV2 U4 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV2 U5 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U7 ( .I(n9), .ZN(n2) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_85 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_85 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_613 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_612 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_611 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_610 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_609 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_608 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_607 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_84 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_606 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_605 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_604 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_XOR2HSV0 U1 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U2 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U5 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0SR U6 ( .I(n8), .ZN(n4) );
  LVT_INHSV2 U7 ( .I(t_i_1_in), .ZN(n5) );
  LVT_CLKNAND2HSV1 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_603 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_602 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_601 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_600 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module row_other_84 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_84 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_606 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_605 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_604 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_603 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_602 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_601 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_600 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_12 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_12 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(
        t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), 
        .t_i_1_out(t0), .t_i_2_out(t_i_2_out[6]) );
  row_other_90 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_89 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_88 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_87 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_86 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_85 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_84 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_73 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_72 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_7bit_48 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module PE_12 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, 
        t_i_2_in, a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro
 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  regist_8bit_77 u0 ( .clk(clk), .rstn(n18), .in(a_in), .out(l_a) );
  regist_8bit_76 u1 ( .clk(clk), .rstn(n18), .in(b_in), .out(b_out) );
  regist_8bit_75 u2 ( .clk(clk), .rstn(n18), .in(g_in), .out(l_g) );
  regist_1bit_51 u3 ( .clk(clk), .rstn(n18), .in(ctr), .out(l_ctr) );
  regist_1bit_50 u4 ( .clk(clk), .rstn(n18), .in(n15), .out(ctro) );
  regist_7bit_51 u5 ( .clk(clk), .rstn(n18), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_7bit_50 u6 ( .clk(clk), .rstn(n18), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_49 u7 ( .clk(clk), .rstn(n18), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_8bit_74 u9 ( .clk(clk), .rstn(n18), .in(mux_b), .out(mux_bq) );
  regist_1bit_48 u10 ( .clk(clk), .rstn(n18), .in(n14), .out(ti_1) );
  regist_7bit_49 u11 ( .clk(clk), .rstn(n18), .in(to_7), .out(ti_7) );
  PE_core_12 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out(t_i_2_out), .t_i_1_out_0(t_i_1_out_0)
         );
  regist_8bit_73 u12 ( .clk(clk), .rstn(n18), .in(ao), .out(a_out) );
  regist_8bit_72 u13 ( .clk(clk), .rstn(n18), .in(go), .out(g_out) );
  regist_7bit_48 u14 ( .clk(clk), .rstn(n18), .in(to), .out(t_i_1_out) );
  LVT_CLKNAND2HSV4 U2 ( .A1(t_i_2_out[0]), .A2(n24), .ZN(n17) );
  LVT_NAND2HSV2 U3 ( .A1(ti_7[1]), .A2(ctro), .ZN(n10) );
  LVT_NAND2HSV8 U4 ( .A1(n10), .A2(n11), .ZN(to_7[1]) );
  LVT_NOR3HSV2 U5 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), 
        .ZN(n21) );
  LVT_AOI21HSV2 U6 ( .A1(n20), .A2(n21), .B(n22), .ZN(\c_t_i_1_in[0] ) );
  LVT_NAND2HSV2 U7 ( .A1(ti_7[0]), .A2(ctro), .ZN(n16) );
  LVT_NAND2HSV2 U8 ( .A1(t_i_2_out[5]), .A2(n24), .ZN(n9) );
  LVT_INHSV2 U9 ( .I(ctro), .ZN(n24) );
  LVT_NAND2HSV8 U10 ( .A1(n17), .A2(n16), .ZN(to_7[0]) );
  LVT_CLKNAND2HSV1 U11 ( .A1(ti_7[3]), .A2(ctro), .ZN(n6) );
  LVT_CLKNAND2HSV3 U12 ( .A1(t_i_2_out[3]), .A2(n24), .ZN(n7) );
  LVT_NAND2HSV4 U13 ( .A1(n6), .A2(n7), .ZN(to_7[3]) );
  LVT_NAND2HSV0P5 U14 ( .A1(ti_7[5]), .A2(ctro), .ZN(n8) );
  LVT_NAND2HSV4 U15 ( .A1(n8), .A2(n9), .ZN(to_7[5]) );
  LVT_NAND2HSV4 U16 ( .A1(t_i_2_out[1]), .A2(n24), .ZN(n11) );
  LVT_INHSV4 U17 ( .I(l_t_i_1_in_0), .ZN(n23) );
  LVT_NOR4HSV12 U18 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(
        l_t_i_1_in[4]), .A4(l_t_i_1_in[3]), .ZN(n20) );
  LVT_INHSV6 U19 ( .I(n19), .ZN(n18) );
  LVT_BUFHSV2RT U20 ( .I(n22), .Z(n12) );
  LVT_INHSV0SR U21 ( .I(l_ctr), .ZN(n22) );
  LVT_INHSV0SR U22 ( .I(to_1), .ZN(n13) );
  LVT_INHSV2 U23 ( .I(n13), .ZN(n14) );
  LVT_AO22HSV1 U24 ( .A1(mux_bq[0]), .A2(n15), .B1(b_out[0]), .B2(n12), .Z(
        mux_b[0]) );
  LVT_AO22HSV1 U25 ( .A1(mux_bq[4]), .A2(n15), .B1(b_out[4]), .B2(n12), .Z(
        mux_b[4]) );
  LVT_AO22HSV1 U26 ( .A1(mux_bq[3]), .A2(n15), .B1(b_out[3]), .B2(n12), .Z(
        mux_b[3]) );
  LVT_AO22HSV1 U27 ( .A1(mux_bq[2]), .A2(n15), .B1(b_out[2]), .B2(n12), .Z(
        mux_b[2]) );
  LVT_AO22HSV1 U28 ( .A1(mux_bq[1]), .A2(n15), .B1(b_out[1]), .B2(n12), .Z(
        mux_b[1]) );
  LVT_AO22HSV1 U29 ( .A1(mux_bq[7]), .A2(n15), .B1(b_out[7]), .B2(n12), .Z(
        mux_b[7]) );
  LVT_AO22HSV1 U30 ( .A1(mux_bq[6]), .A2(n15), .B1(b_out[6]), .B2(n12), .Z(
        mux_b[6]) );
  LVT_AO22HSV1 U31 ( .A1(mux_bq[5]), .A2(n15), .B1(b_out[5]), .B2(n12), .Z(
        mux_b[5]) );
  LVT_NOR2HSV0 U32 ( .A1(n23), .A2(n22), .ZN(c_t_i_1_in_0) );
  LVT_MOAI22HSV4 U33 ( .A1(l_ctr), .A2(n23), .B1(ti_1), .B2(l_ctr), .ZN(to_1)
         );
  LVT_INHSV2 U34 ( .I(n22), .ZN(n15) );
  LVT_AO22HSV4 U35 ( .A1(ti_7[2]), .A2(ctro), .B1(t_i_2_out[2]), .B2(n24), .Z(
        to_7[2]) );
  LVT_AO22HSV4 U36 ( .A1(ti_7[4]), .A2(ctro), .B1(t_i_2_out[4]), .B2(n24), .Z(
        to_7[4]) );
  LVT_AO22HSV4 U37 ( .A1(ti_7[6]), .A2(ctro), .B1(t_i_2_out[6]), .B2(n24), .Z(
        to_7[6]) );
  LVT_INHSV2 U38 ( .I(rstn), .ZN(n19) );
endmodule


module regist_8bit_71 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_70 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_69 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_47 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_46 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV1 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_47 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_46 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
endmodule


module regist_1bit_45 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_68 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_44 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_45 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module cell_3_599 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_83 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_82 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n2), .A3(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_81 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U3 ( .A1(n5), .A2(n6), .Z(n7) );
endmodule


module cell_4_80 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_79 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_XOR3HSV1 U2 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
endmodule


module cell_4_78 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_XOR3HSV1 U2 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
endmodule


module cell_4_77 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n7), .A2(n1), .ZN(t_i_out) );
  LVT_CLKXOR2HSV4 U3 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_XNOR2HSV1 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n1) );
endmodule


module row_1_11 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_3_599 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_83 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(
        t_i_1_out[1]) );
  cell_4_82 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_81 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(
        t_i_1_out[3]) );
  cell_4_80 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(
        t_i_1_out[4]) );
  cell_4_79 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(t_i_1_out[5])
         );
  cell_4_78 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_77 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_CLKNHSV0P5 U2 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U3 ( .I(n2), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n4) );
endmodule


module cell_2_83 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_598 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_597 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_596 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_595 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_594 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_593 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV1 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_592 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_CLKNAND2HSV1 U1 ( .A1(n4), .A2(n5), .ZN(t_i_out) );
  LVT_INAND2HSV2 U2 ( .A1(n6), .B1(n2), .ZN(n5) );
  LVT_INHSV4SR U4 ( .I(n8), .ZN(n2) );
  LVT_CLKNAND2HSV3 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U6 ( .A1(n6), .A2(n8), .ZN(n4) );
  LVT_XNOR2HSV4 U7 ( .A1(t_i_1_in), .A2(n7), .ZN(n6) );
endmodule


module row_other_83 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_83 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_598 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_597 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_596 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_595 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_594 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_593 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_592 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_82 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_591 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_590 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_589 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_588 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_587 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XOR2HSV0 U4 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_586 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_585 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKNAND2HSV2 U2 ( .A1(n5), .A2(n4), .ZN(t_i_out) );
  LVT_INAND2HSV2 U4 ( .A1(n8), .B1(n2), .ZN(n5) );
  LVT_INHSV2 U5 ( .I(n6), .ZN(n2) );
  LVT_CLKNAND2HSV1 U6 ( .A1(n6), .A2(n8), .ZN(n4) );
  LVT_XNOR2HSV4 U7 ( .A1(t_i_1_in), .A2(n7), .ZN(n6) );
endmodule


module row_other_82 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_82 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_591 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_590 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_589 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_588 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_587 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_586 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_585 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_81 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_584 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_583 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_582 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_581 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_580 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_579 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_OAI21HSV2 U1 ( .A1(t_i_1_in), .A2(n5), .B(n2), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_NAND2HSV0 U4 ( .A1(n5), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV4 U5 ( .A1(n6), .A2(n4), .ZN(t_i_out) );
endmodule


module cell_3_578 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_IOA21HSV4 U2 ( .A1(n8), .A2(n6), .B(n5), .ZN(t_i_out) );
  LVT_INHSV2P5 U4 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV4 U5 ( .A1(n2), .A2(n4), .ZN(n5) );
  LVT_XNOR2HSV4 U6 ( .A1(t_i_1_in), .A2(n7), .ZN(n6) );
  LVT_INHSV3SR U7 ( .I(n8), .ZN(n2) );
endmodule


module row_other_81 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_81 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_584 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_583 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_582 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_581 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_580 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_579 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_578 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_80 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_577 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_576 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_575 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_574 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_573 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_572 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_571 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_NAND2HSV4 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module row_other_80 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_80 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_577 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_576 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_575 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_574 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_573 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_572 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_571 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_79 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_570 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_569 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKXOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_568 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_567 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_566 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_565 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XNOR2HSV4 U2 ( .A1(n6), .A2(n4), .ZN(t_i_out) );
  LVT_OAI21HSV2 U4 ( .A1(t_i_1_in), .A2(n5), .B(n2), .ZN(n4) );
  LVT_NAND2HSV2 U5 ( .A1(n5), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_564 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV3SR U2 ( .I(n9), .ZN(n2) );
  LVT_INHSV3SR U4 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV4 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV4 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U7 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNAND2HSV3 U8 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
endmodule


module row_other_79 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_79 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_570 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_569 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_568 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_567 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_566 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_565 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_564 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_78 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_563 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_562 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_561 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_560 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_559 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_558 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_557 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module row_other_78 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_78 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_563 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_562 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_561 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_560 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_559 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_558 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_557 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_77 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_556 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n8), .Z(n9) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV0P5 U4 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_NAND2HSV1 U6 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV0P5SR U7 ( .I(n10), .ZN(n4) );
  LVT_INHSV0SR U8 ( .I(n9), .ZN(n5) );
endmodule


module cell_3_555 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_554 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_553 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_552 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_551 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKXOR2HSV2 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_550 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module row_other_77 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_77 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_556 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_555 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_554 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_553 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_552 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_551 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_550 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_11 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_11 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(
        t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), 
        .t_i_1_out(t0), .t_i_2_out(t_i_2_out[6]) );
  row_other_83 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_82 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_81 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_80 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_79 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_78 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_77 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_67 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_66 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_7bit_44 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module PE_11 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, 
        t_i_2_in, a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro
 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  regist_8bit_71 u0 ( .clk(clk), .rstn(n17), .in(a_in), .out(l_a) );
  regist_8bit_70 u1 ( .clk(clk), .rstn(n17), .in(b_in), .out(b_out) );
  regist_8bit_69 u2 ( .clk(clk), .rstn(n17), .in(g_in), .out(l_g) );
  regist_1bit_47 u3 ( .clk(clk), .rstn(n17), .in(ctr), .out(l_ctr) );
  regist_1bit_46 u4 ( .clk(clk), .rstn(n17), .in(n14), .out(ctro) );
  regist_7bit_47 u5 ( .clk(clk), .rstn(n17), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_7bit_46 u6 ( .clk(clk), .rstn(n17), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_45 u7 ( .clk(clk), .rstn(n17), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_8bit_68 u9 ( .clk(clk), .rstn(n17), .in(mux_b), .out(mux_bq) );
  regist_1bit_44 u10 ( .clk(clk), .rstn(n17), .in(to_1), .out(ti_1) );
  regist_7bit_45 u11 ( .clk(clk), .rstn(n17), .in(to_7), .out(ti_7) );
  PE_core_11 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out(t_i_2_out), .t_i_1_out_0(t_i_1_out_0)
         );
  regist_8bit_67 u12 ( .clk(clk), .rstn(n17), .in(ao), .out(a_out) );
  regist_8bit_66 u13 ( .clk(clk), .rstn(n17), .in(go), .out(g_out) );
  regist_7bit_44 u14 ( .clk(clk), .rstn(n17), .in(to), .out(t_i_1_out) );
  LVT_INHSV4SR U2 ( .I(l_t_i_1_in_0), .ZN(n22) );
  LVT_INHSV4 U3 ( .I(n12), .ZN(n13) );
  LVT_INHSV2 U4 ( .I(n21), .ZN(n12) );
  LVT_NAND2HSV2 U5 ( .A1(ti_7[0]), .A2(ctro), .ZN(n15) );
  LVT_NAND2HSV4 U6 ( .A1(t_i_2_out[0]), .A2(n23), .ZN(n16) );
  LVT_NAND2HSV8 U7 ( .A1(n16), .A2(n15), .ZN(to_7[0]) );
  LVT_NAND2HSV8 U8 ( .A1(n10), .A2(n11), .ZN(to_7[6]) );
  LVT_NAND2HSV8 U9 ( .A1(n6), .A2(n7), .ZN(to_7[4]) );
  LVT_NOR4HSV12 U10 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(
        l_t_i_1_in[4]), .A4(l_t_i_1_in[3]), .ZN(n19) );
  LVT_INHSV2 U11 ( .I(ctro), .ZN(n23) );
  LVT_NAND2HSV4 U12 ( .A1(t_i_2_out[4]), .A2(n23), .ZN(n7) );
  LVT_NAND2HSV2 U13 ( .A1(ti_7[4]), .A2(ctro), .ZN(n6) );
  LVT_NOR2HSV2 U14 ( .A1(l_t_i_1_in[1]), .A2(l_t_i_1_in[2]), .ZN(n8) );
  LVT_NOR2HSV2 U15 ( .A1(l_t_i_1_in[0]), .A2(n9), .ZN(n20) );
  LVT_INHSV2 U16 ( .I(n8), .ZN(n9) );
  LVT_AOI21HSV2 U17 ( .A1(n20), .A2(n19), .B(n13), .ZN(\c_t_i_1_in[0] ) );
  LVT_NAND2HSV2 U18 ( .A1(ti_7[6]), .A2(ctro), .ZN(n10) );
  LVT_CLKNAND2HSV4 U19 ( .A1(t_i_2_out[6]), .A2(n23), .ZN(n11) );
  LVT_INHSV6 U20 ( .I(n18), .ZN(n17) );
  LVT_NOR2HSV0 U21 ( .A1(n22), .A2(n13), .ZN(c_t_i_1_in_0) );
  LVT_CLKNHSV1 U22 ( .I(l_ctr), .ZN(n21) );
  LVT_CLKNHSV1 U23 ( .I(n13), .ZN(n14) );
  LVT_AO22HSV2 U24 ( .A1(mux_bq[4]), .A2(n14), .B1(b_out[4]), .B2(n13), .Z(
        mux_b[4]) );
  LVT_AO22HSV2 U25 ( .A1(mux_bq[1]), .A2(n14), .B1(b_out[1]), .B2(n13), .Z(
        mux_b[1]) );
  LVT_AO22HSV2 U26 ( .A1(mux_bq[0]), .A2(n14), .B1(b_out[0]), .B2(n13), .Z(
        mux_b[0]) );
  LVT_AO22HSV2 U27 ( .A1(mux_bq[7]), .A2(l_ctr), .B1(b_out[7]), .B2(n13), .Z(
        mux_b[7]) );
  LVT_AO22HSV2 U28 ( .A1(mux_bq[6]), .A2(l_ctr), .B1(b_out[6]), .B2(n13), .Z(
        mux_b[6]) );
  LVT_AO22HSV2 U29 ( .A1(mux_bq[5]), .A2(l_ctr), .B1(b_out[5]), .B2(n13), .Z(
        mux_b[5]) );
  LVT_AO22HSV2 U30 ( .A1(mux_bq[3]), .A2(n14), .B1(b_out[3]), .B2(n13), .Z(
        mux_b[3]) );
  LVT_AO22HSV2 U31 ( .A1(mux_bq[2]), .A2(n14), .B1(b_out[2]), .B2(n13), .Z(
        mux_b[2]) );
  LVT_AO22HSV4 U32 ( .A1(ti_7[1]), .A2(ctro), .B1(t_i_2_out[1]), .B2(n23), .Z(
        to_7[1]) );
  LVT_AO22HSV4 U33 ( .A1(ti_7[2]), .A2(ctro), .B1(t_i_2_out[2]), .B2(n23), .Z(
        to_7[2]) );
  LVT_AO22HSV4 U34 ( .A1(ti_7[3]), .A2(ctro), .B1(t_i_2_out[3]), .B2(n23), .Z(
        to_7[3]) );
  LVT_AO22HSV4 U35 ( .A1(ti_7[5]), .A2(ctro), .B1(t_i_2_out[5]), .B2(n23), .Z(
        to_7[5]) );
  LVT_MOAI22HSV4 U36 ( .A1(l_ctr), .A2(n22), .B1(ti_1), .B2(l_ctr), .ZN(to_1)
         );
  LVT_INHSV2 U37 ( .I(rstn), .ZN(n18) );
endmodule


module regist_8bit_65 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_64 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_63 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_43 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_42 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_43 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV4 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_42 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
endmodule


module regist_1bit_41 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_62 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_40 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_41 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module cell_3_549 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_76 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U3 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_75 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_74 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_73 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_72 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_71 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n9) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n8), .A2(n9), .Z(n10) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_INAND2HSV2 U3 ( .A1(n7), .B1(n1), .ZN(n6) );
  LVT_NAND2HSV2 U5 ( .A1(n7), .A2(n10), .ZN(n5) );
  LVT_NAND2HSV2 U6 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV2 U7 ( .I(n10), .ZN(n1) );
  LVT_XNOR2HSV1 U8 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n7) );
endmodule


module cell_4_70 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10, n11;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n10) );
  LVT_CLKNHSV1 U1 ( .I(n9), .ZN(n6) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV4 U3 ( .A1(n11), .A2(n1), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n1) );
  LVT_NAND2HSV0P5 U6 ( .A1(n10), .A2(n6), .ZN(n7) );
  LVT_NAND2HSV0 U7 ( .A1(n5), .A2(n9), .ZN(n8) );
  LVT_NAND2HSV2 U8 ( .A1(n7), .A2(n8), .ZN(n11) );
  LVT_INHSV0SR U9 ( .I(n10), .ZN(n5) );
endmodule


module row_1_10 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_3_549 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_76 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(
        t_i_1_out[1]) );
  cell_4_75 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_74 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(
        t_i_1_out[3]) );
  cell_4_73 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(
        t_i_1_out[4]) );
  cell_4_72 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(
        t_i_1_out[5]) );
  cell_4_71 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_70 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_76 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_548 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_547 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_546 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_545 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_544 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_543 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_542 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4;

  LVT_XOR2HSV2 U1 ( .A1(n2), .A2(t_i_1_in), .Z(n3) );
  LVT_NAND2HSV3 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n4) );
  LVT_CLKAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .Z(n2) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(n3), .ZN(t_i_out) );
endmodule


module row_other_76 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_76 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_548 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_547 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_546 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_545 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_544 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_543 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_542 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_75 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_541 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_540 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_539 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_538 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_537 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_536 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_INHSV2 U1 ( .I(t_i_1_in), .ZN(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n9), .A2(n10), .Z(t_i_out) );
  LVT_NAND2HSV2 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV0P5 U4 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U6 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV2 U7 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0 U8 ( .A1(b_in), .A2(a_in), .ZN(n8) );
endmodule


module cell_3_535 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U1 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV4 U5 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV3SR U6 ( .I(n9), .ZN(n2) );
  LVT_INHSV4SR U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_75 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_75 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_541 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_540 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_539 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_538 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_537 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_536 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_535 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_74 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_534 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_533 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_532 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_531 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_530 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_529 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_528 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV4 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV1 U5 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
  LVT_NAND2HSV2 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U7 ( .I(n9), .ZN(n2) );
  LVT_INHSV2 U8 ( .I(n7), .ZN(n4) );
endmodule


module row_other_74 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_74 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_534 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_533 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_532 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_531 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_530 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_529 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_528 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_73 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_527 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_526 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_525 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_524 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_523 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_522 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKXOR2HSV2 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_521 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNHSV2P5 U1 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV4 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV0P5 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV3SR U5 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV4 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_73 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_73 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_527 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_526 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_525 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_524 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_523 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_522 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_521 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_72 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_520 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_519 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_518 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_517 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_516 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_515 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_514 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4, n5, n6, n7, n8;

  LVT_INHSV2SR U1 ( .I(n8), .ZN(n2) );
  LVT_NAND2HSV0P5 U2 ( .A1(n8), .A2(n6), .ZN(n4) );
  LVT_NAND2HSV2 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_INHSV2 U4 ( .I(n6), .ZN(n3) );
  LVT_NAND2HSV4 U5 ( .A1(n4), .A2(n5), .ZN(t_i_out) );
  LVT_CLKAND2HSV2 U6 ( .A1(b_in), .A2(a_in), .Z(n7) );
  LVT_CLKXOR2HSV4 U7 ( .A1(t_i_1_in), .A2(n7), .Z(n6) );
  LVT_NAND2HSV4 U8 ( .A1(n2), .A2(n3), .ZN(n5) );
endmodule


module row_other_72 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_72 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_520 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_519 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_518 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_517 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_516 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_515 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_514 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_71 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_513 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_512 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_511 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_510 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_509 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_508 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_507 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U5 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV0P5 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2SR U7 ( .I(n9), .ZN(n2) );
  LVT_INHSV2 U8 ( .I(n7), .ZN(n4) );
endmodule


module row_other_71 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_71 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_513 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_512 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_511 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_510 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_509 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_508 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_507 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_70 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_506 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_505 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_504 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_503 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_502 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_501 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_500 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module row_other_70 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_70 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_506 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_505 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_504 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_503 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_502 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_501 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_500 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_10 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_10 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(
        t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), 
        .t_i_1_out(t0), .t_i_2_out(t_i_2_out[6]) );
  row_other_76 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_75 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_74 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_73 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_72 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_71 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_70 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_61 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_60 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_7bit_40 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
endmodule


module PE_10 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, 
        t_i_2_in, a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro
 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  LVT_NOR3HSV0 U24 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), .ZN(n17) );
  regist_8bit_65 u0 ( .clk(clk), .rstn(n14), .in(a_in), .out(l_a) );
  regist_8bit_64 u1 ( .clk(clk), .rstn(n14), .in(b_in), .out(b_out) );
  regist_8bit_63 u2 ( .clk(clk), .rstn(n14), .in(g_in), .out(l_g) );
  regist_1bit_43 u3 ( .clk(clk), .rstn(n14), .in(ctr), .out(l_ctr) );
  regist_1bit_42 u4 ( .clk(clk), .rstn(n14), .in(n11), .out(ctro) );
  regist_7bit_43 u5 ( .clk(clk), .rstn(n14), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_7bit_42 u6 ( .clk(clk), .rstn(n14), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_41 u7 ( .clk(clk), .rstn(n14), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_8bit_62 u9 ( .clk(clk), .rstn(n14), .in(mux_b), .out(mux_bq) );
  regist_1bit_40 u10 ( .clk(clk), .rstn(n14), .in(n9), .out(ti_1) );
  regist_7bit_41 u11 ( .clk(clk), .rstn(n14), .in(to_7), .out(ti_7) );
  PE_core_10 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out(t_i_2_out), .t_i_1_out_0(t_i_1_out_0)
         );
  regist_8bit_61 u12 ( .clk(clk), .rstn(n14), .in(ao), .out(a_out) );
  regist_8bit_60 u13 ( .clk(clk), .rstn(n14), .in(go), .out(g_out) );
  regist_7bit_40 u14 ( .clk(clk), .rstn(n14), .in(to), .out(t_i_1_out) );
  LVT_NAND2HSV2 U2 ( .A1(ti_7[1]), .A2(ctro), .ZN(n6) );
  LVT_CLKNAND2HSV4 U3 ( .A1(t_i_2_out[1]), .A2(n20), .ZN(n7) );
  LVT_INHSV2 U4 ( .I(ctro), .ZN(n20) );
  LVT_NOR4HSV12 U5 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(l_t_i_1_in[4]), .A4(l_t_i_1_in[3]), .ZN(n16) );
  LVT_NAND2HSV8 U6 ( .A1(n7), .A2(n6), .ZN(to_7[1]) );
  LVT_NAND2HSV2 U7 ( .A1(ti_7[5]), .A2(ctro), .ZN(n12) );
  LVT_NAND2HSV4 U8 ( .A1(t_i_2_out[5]), .A2(n20), .ZN(n13) );
  LVT_INHSV6 U9 ( .I(n15), .ZN(n14) );
  LVT_INHSV0SR U10 ( .I(to_1), .ZN(n8) );
  LVT_INHSV2 U11 ( .I(n8), .ZN(n9) );
  LVT_BUFHSV2RT U12 ( .I(n18), .Z(n10) );
  LVT_INHSV0SR U13 ( .I(l_ctr), .ZN(n18) );
  LVT_NOR2HSV2 U14 ( .A1(n19), .A2(n18), .ZN(c_t_i_1_in_0) );
  LVT_AOI21HSV1 U15 ( .A1(n17), .A2(n16), .B(n18), .ZN(\c_t_i_1_in[0] ) );
  LVT_MOAI22HSV4 U16 ( .A1(l_ctr), .A2(n19), .B1(ti_1), .B2(l_ctr), .ZN(to_1)
         );
  LVT_CLKNAND2HSV8 U17 ( .A1(n13), .A2(n12), .ZN(to_7[5]) );
  LVT_INHSV3SR U18 ( .I(l_t_i_1_in_0), .ZN(n19) );
  LVT_INHSV2 U19 ( .I(n18), .ZN(n11) );
  LVT_AO22HSV2 U20 ( .A1(mux_bq[0]), .A2(n11), .B1(b_out[0]), .B2(n10), .Z(
        mux_b[0]) );
  LVT_AO22HSV2 U21 ( .A1(mux_bq[1]), .A2(n11), .B1(b_out[1]), .B2(n10), .Z(
        mux_b[1]) );
  LVT_AO22HSV2 U22 ( .A1(mux_bq[2]), .A2(n11), .B1(b_out[2]), .B2(n10), .Z(
        mux_b[2]) );
  LVT_AO22HSV2 U23 ( .A1(mux_bq[3]), .A2(n11), .B1(b_out[3]), .B2(n10), .Z(
        mux_b[3]) );
  LVT_AO22HSV2 U25 ( .A1(mux_bq[4]), .A2(n11), .B1(b_out[4]), .B2(n10), .Z(
        mux_b[4]) );
  LVT_AO22HSV2 U26 ( .A1(mux_bq[5]), .A2(n11), .B1(b_out[5]), .B2(n10), .Z(
        mux_b[5]) );
  LVT_AO22HSV2 U27 ( .A1(mux_bq[6]), .A2(n11), .B1(b_out[6]), .B2(n10), .Z(
        mux_b[6]) );
  LVT_AO22HSV2 U28 ( .A1(mux_bq[7]), .A2(n11), .B1(b_out[7]), .B2(n18), .Z(
        mux_b[7]) );
  LVT_AO22HSV4 U29 ( .A1(ti_7[0]), .A2(ctro), .B1(t_i_2_out[0]), .B2(n20), .Z(
        to_7[0]) );
  LVT_AO22HSV4 U30 ( .A1(ti_7[2]), .A2(ctro), .B1(t_i_2_out[2]), .B2(n20), .Z(
        to_7[2]) );
  LVT_AO22HSV4 U31 ( .A1(ti_7[3]), .A2(ctro), .B1(t_i_2_out[3]), .B2(n20), .Z(
        to_7[3]) );
  LVT_AO22HSV4 U32 ( .A1(ti_7[4]), .A2(ctro), .B1(t_i_2_out[4]), .B2(n20), .Z(
        to_7[4]) );
  LVT_AO22HSV4 U33 ( .A1(ti_7[6]), .A2(ctro), .B1(t_i_2_out[6]), .B2(n20), .Z(
        to_7[6]) );
  LVT_INHSV2 U34 ( .I(rstn), .ZN(n15) );
endmodule


module regist_8bit_59 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_58 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_57 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_39 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_38 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_39 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_38 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
endmodule


module regist_1bit_37 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_56 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_36 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_37 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module cell_3_499 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_69 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_XOR2HSV2 U2 ( .A1(t_i_1_in), .A2(t_i_2_in), .Z(n8) );
  LVT_XOR2HSV2 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_68 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_67 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_66 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV2 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_65 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV4 U1 ( .A1(n7), .A2(n8), .Z(t_i_out) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_64 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U3 ( .A1(n1), .A2(n7), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n1) );
endmodule


module cell_4_63 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10, n11;

  LVT_CLKNHSV2 U1 ( .I(n9), .ZN(n1) );
  LVT_CLKNAND2HSV3 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV3 U3 ( .A1(n7), .A2(n6), .ZN(n11) );
  LVT_NAND2HSV0P5 U4 ( .A1(n5), .A2(n9), .ZN(n6) );
  LVT_NAND2HSV2 U5 ( .A1(b_in), .A2(a_in), .ZN(n10) );
  LVT_CLKNAND2HSV2 U6 ( .A1(n1), .A2(n10), .ZN(n7) );
  LVT_INHSV0SR U7 ( .I(n10), .ZN(n5) );
  LVT_XNOR2HSV4 U8 ( .A1(n11), .A2(n8), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U9 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n8) );
endmodule


module row_1_9 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_3_499 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_69 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(
        t_i_1_out[1]) );
  cell_4_68 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_67 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(
        t_i_1_out[3]) );
  cell_4_66 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(
        t_i_1_out[4]) );
  cell_4_65 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(
        t_i_1_out[5]) );
  cell_4_64 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_63 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_69 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_498 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_497 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_496 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_495 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_494 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_493 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_492 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4, n5, n6, n7, n8;

  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_INHSV2SR U2 ( .I(n8), .ZN(n2) );
  LVT_CLKNAND2HSV3 U3 ( .A1(n4), .A2(n5), .ZN(t_i_out) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n6), .Z(n7) );
  LVT_INHSV2 U5 ( .I(n7), .ZN(n3) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n2), .A2(n3), .ZN(n5) );
  LVT_AND2HSV0RD U7 ( .A1(b_in), .A2(a_in), .Z(n6) );
  LVT_NAND2HSV0P5 U8 ( .A1(n8), .A2(n7), .ZN(n4) );
endmodule


module row_other_69 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_69 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_498 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_497 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_496 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_495 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_494 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_493 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_492 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_68 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_491 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_490 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_489 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_488 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_487 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_486 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_485 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_INHSV3SR U4 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV4SR U6 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U7 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV4 U8 ( .A1(n2), .A2(n4), .ZN(n6) );
endmodule


module row_other_68 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_68 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_491 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_490 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_489 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_488 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_487 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_486 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_485 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_67 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_484 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_483 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_482 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_481 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_480 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_479 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_478 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV4 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV2 U2 ( .I(n7), .ZN(n4) );
  LVT_INHSV4SR U4 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV4 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV0P5 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV4 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_67 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_67 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_484 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_483 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_482 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_481 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_480 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_479 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_478 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV2 U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV0P5SR U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_66 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_477 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_476 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_475 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_474 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_473 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_472 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_471 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U1 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV2 U4 ( .I(n9), .ZN(n2) );
  LVT_CLKNHSV2 U5 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV4 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_66 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_66 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_477 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_476 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_475 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_474 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_473 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_472 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_471 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_65 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_470 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV1 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_469 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_468 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_467 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_466 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_465 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_464 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U1 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV4SR U2 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV2 U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV4 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV4 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_65 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_65 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_470 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_469 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_468 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_467 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_466 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_465 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_464 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_64 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n1, n3;

  LVT_XNOR2HSV4 U1 ( .A1(n3), .A2(n1), .ZN(t_i_out) );
  LVT_CLKAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .Z(n1) );
  LVT_CLKNAND2HSV0 U3 ( .A1(g_in), .A2(t_m_1_in), .ZN(n3) );
endmodule


module cell_3_463 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_462 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_461 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_460 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_459 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_458 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_457 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV2 U1 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV4SR U5 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV4 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV4 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_64 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_64 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_463 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_462 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_461 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_460 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_459 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_458 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_457 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_63 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n1, n3;

  LVT_XNOR2HSV1 U1 ( .A1(n3), .A2(n1), .ZN(t_i_out) );
  LVT_AND2HSV32 U2 ( .A1(b_in), .A2(a_in), .Z(n1) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_456 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_455 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNHSV2 U1 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_CLKNAND2HSV1 U4 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_XOR2HSV2 U5 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_CLKNHSV0 U6 ( .I(n10), .ZN(n4) );
  LVT_NAND2HSV2 U7 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U8 ( .A1(n10), .A2(n5), .ZN(n6) );
endmodule


module cell_3_454 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module cell_3_453 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9;

  LVT_XOR2HSV0 U1 ( .A1(n9), .A2(n8), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_INAND2HSV2 U2 ( .A1(t_i_1_in), .B1(n7), .ZN(n6) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U5 ( .A1(t_i_1_in), .A2(n4), .ZN(n5) );
  LVT_NAND2HSV2 U6 ( .A1(n5), .A2(n6), .ZN(n8) );
  LVT_INHSV2 U7 ( .I(n7), .ZN(n4) );
endmodule


module cell_3_452 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_451 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV1 U2 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV2 U4 ( .I(n9), .ZN(n5) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_INHSV0P5SR U6 ( .I(n10), .ZN(n4) );
  LVT_NAND2HSV0P5 U7 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_XOR2HSV2 U8 ( .A1(t_i_1_in), .A2(n8), .Z(n9) );
endmodule


module cell_3_450 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKXOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module row_other_63 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_63 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_456 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_455 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_454 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_453 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_452 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_451 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_450 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_9 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_9 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), .t_i_1_out(t0), 
        .t_i_2_out(t_i_2_out[6]) );
  row_other_69 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_68 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_67 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_66 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_65 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_64 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_63 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_55 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_54 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_7bit_36 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module PE_9 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   n23, n24, l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1,
         ti_1, n2, n6, n7, n8, n9, n10, n11, n12, n13, n15, n17, n18, n19, n20,
         n21, n22;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  LVT_NOR3HSV0 U24 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), .ZN(n20) );
  regist_8bit_59 u0 ( .clk(clk), .rstn(n17), .in(a_in), .out(l_a) );
  regist_8bit_58 u1 ( .clk(clk), .rstn(n17), .in(b_in), .out(b_out) );
  regist_8bit_57 u2 ( .clk(clk), .rstn(n17), .in(g_in), .out(l_g) );
  regist_1bit_39 u3 ( .clk(clk), .rstn(n17), .in(ctr), .out(l_ctr) );
  regist_1bit_38 u4 ( .clk(clk), .rstn(n17), .in(n12), .out(ctro) );
  regist_7bit_39 u5 ( .clk(clk), .rstn(n17), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_7bit_38 u6 ( .clk(clk), .rstn(n17), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_37 u7 ( .clk(clk), .rstn(n17), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_8bit_56 u9 ( .clk(clk), .rstn(n17), .in(mux_b), .out(mux_bq) );
  regist_1bit_36 u10 ( .clk(clk), .rstn(n17), .in(n11), .out(ti_1) );
  regist_7bit_37 u11 ( .clk(clk), .rstn(n17), .in(to_7), .out(ti_7) );
  PE_core_9 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out({t_i_2_out[6], n23, t_i_2_out[4:3], 
        n24, t_i_2_out[1:0]}), .t_i_1_out_0(t_i_1_out_0) );
  regist_8bit_55 u12 ( .clk(clk), .rstn(n17), .in(ao), .out(a_out) );
  regist_8bit_54 u13 ( .clk(clk), .rstn(n17), .in(go), .out(g_out) );
  regist_7bit_36 u14 ( .clk(clk), .rstn(n17), .in(to), .out(t_i_1_out) );
  LVT_NAND2HSV8 U2 ( .A1(t_i_2_out[3]), .A2(n22), .ZN(n7) );
  LVT_IOA22HSV4 U3 ( .B1(l_ctr), .B2(n10), .A1(ti_1), .A2(l_ctr), .ZN(to_1) );
  LVT_NOR4HSV12 U4 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(l_t_i_1_in[4]), .A4(l_t_i_1_in[3]), .ZN(n19) );
  LVT_INHSV2 U5 ( .I(n8), .ZN(n2) );
  LVT_AOI21HSV2 U6 ( .A1(n20), .A2(n19), .B(n9), .ZN(\c_t_i_1_in[0] ) );
  LVT_BUFHSV2 U7 ( .I(n21), .Z(n8) );
  LVT_INHSV2 U8 ( .I(ctro), .ZN(n22) );
  LVT_AO22HSV1 U9 ( .A1(mux_bq[5]), .A2(n2), .B1(b_out[5]), .B2(n9), .Z(
        mux_b[5]) );
  LVT_NAND2HSV4 U10 ( .A1(ti_7[3]), .A2(ctro), .ZN(n6) );
  LVT_NAND2HSV8 U11 ( .A1(n6), .A2(n7), .ZN(to_7[3]) );
  LVT_INHSV4SR U12 ( .I(l_t_i_1_in_0), .ZN(n10) );
  LVT_INHSV6 U13 ( .I(n18), .ZN(n17) );
  LVT_BUFHSV2 U14 ( .I(n21), .Z(n9) );
  LVT_INHSV0SR U15 ( .I(l_ctr), .ZN(n21) );
  LVT_MOAI22HSV0 U16 ( .A1(n2), .A2(n10), .B1(ti_1), .B2(n2), .ZN(n11) );
  LVT_INHSV0SR U17 ( .I(n9), .ZN(n12) );
  LVT_NOR2HSV2 U18 ( .A1(n10), .A2(n8), .ZN(c_t_i_1_in_0) );
  LVT_AO22HSV0 U19 ( .A1(mux_bq[7]), .A2(n12), .B1(b_out[7]), .B2(n9), .Z(
        mux_b[7]) );
  LVT_AO22HSV1 U20 ( .A1(mux_bq[1]), .A2(n12), .B1(b_out[1]), .B2(n8), .Z(
        mux_b[1]) );
  LVT_AO22HSV2 U21 ( .A1(mux_bq[4]), .A2(n12), .B1(b_out[4]), .B2(n8), .Z(
        mux_b[4]) );
  LVT_AO22HSV2 U22 ( .A1(mux_bq[3]), .A2(n12), .B1(b_out[3]), .B2(n8), .Z(
        mux_b[3]) );
  LVT_AO22HSV2 U23 ( .A1(mux_bq[2]), .A2(n12), .B1(b_out[2]), .B2(n8), .Z(
        mux_b[2]) );
  LVT_AO22HSV2 U25 ( .A1(mux_bq[0]), .A2(n12), .B1(b_out[0]), .B2(n8), .Z(
        mux_b[0]) );
  LVT_AO22HSV2 U26 ( .A1(mux_bq[6]), .A2(n2), .B1(b_out[6]), .B2(n9), .Z(
        mux_b[6]) );
  LVT_INHSV0SR U27 ( .I(n24), .ZN(n13) );
  LVT_INHSV2 U28 ( .I(n13), .ZN(t_i_2_out[2]) );
  LVT_INHSV0SR U29 ( .I(n23), .ZN(n15) );
  LVT_INHSV2 U30 ( .I(n15), .ZN(t_i_2_out[5]) );
  LVT_AO22HSV4 U31 ( .A1(ti_7[0]), .A2(ctro), .B1(t_i_2_out[0]), .B2(n22), .Z(
        to_7[0]) );
  LVT_AO22HSV4 U32 ( .A1(ti_7[1]), .A2(ctro), .B1(t_i_2_out[1]), .B2(n22), .Z(
        to_7[1]) );
  LVT_AO22HSV4 U33 ( .A1(ti_7[2]), .A2(ctro), .B1(n24), .B2(n22), .Z(to_7[2])
         );
  LVT_AO22HSV4 U34 ( .A1(ti_7[4]), .A2(ctro), .B1(t_i_2_out[4]), .B2(n22), .Z(
        to_7[4]) );
  LVT_AO22HSV4 U35 ( .A1(ti_7[5]), .A2(ctro), .B1(n23), .B2(n22), .Z(to_7[5])
         );
  LVT_AO22HSV4 U36 ( .A1(ti_7[6]), .A2(ctro), .B1(t_i_2_out[6]), .B2(n22), .Z(
        to_7[6]) );
  LVT_INHSV2 U37 ( .I(rstn), .ZN(n18) );
endmodule


module regist_8bit_53 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_52 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_51 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_35 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_34 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV1 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_35 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_34 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
endmodule


module regist_1bit_33 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_50 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_32 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_33 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module cell_3_449 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_62 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV2 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_61 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_60 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_59 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U3 ( .A1(n6), .A2(n5), .Z(n7) );
endmodule


module cell_4_58 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_57 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n2, n4;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR3HSV1 U1 ( .A1(n1), .A2(n4), .A3(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_XNOR2HSV1 U3 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n1) );
endmodule


module cell_4_56 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  LVT_NAND2HSV2 U1 ( .A1(n10), .A2(n11), .ZN(n15) );
  LVT_NAND2HSV2 U2 ( .A1(n9), .A2(n14), .ZN(n10) );
  LVT_CLKNAND2HSV2 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n13) );
  LVT_CLKNAND2HSV1 U4 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_NAND2HSV2 U5 ( .A1(n1), .A2(n5), .ZN(n7) );
  LVT_NAND2HSV2 U6 ( .A1(b_in), .A2(a_in), .ZN(n14) );
  LVT_XNOR2HSV1 U7 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n12) );
  LVT_INHSV2 U8 ( .I(n15), .ZN(n1) );
  LVT_NAND2HSV1 U9 ( .A1(n15), .A2(n12), .ZN(n6) );
  LVT_INHSV2SR U10 ( .I(n12), .ZN(n5) );
  LVT_CLKNAND2HSV0 U11 ( .A1(n8), .A2(n13), .ZN(n11) );
  LVT_INHSV0SR U12 ( .I(n14), .ZN(n8) );
  LVT_CLKNHSV2 U13 ( .I(n13), .ZN(n9) );
endmodule


module row_1_8 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_3_449 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_62 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(t_i_1_out[1])
         );
  cell_4_61 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_60 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(
        t_i_1_out[3]) );
  cell_4_59 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(
        t_i_1_out[4]) );
  cell_4_58 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(t_i_1_out[5])
         );
  cell_4_57 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(t_i_1_out[6])
         );
  cell_4_56 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
  LVT_INHSV0P5SR U3 ( .I(t_m_1_in), .ZN(n3) );
  LVT_CLKNHSV2 U4 ( .I(n3), .ZN(n4) );
endmodule


module cell_2_62 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_448 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_447 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_446 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_445 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_444 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_443 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_442 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_XNOR2HSV1 U1 ( .A1(t_i_1_in), .A2(n7), .ZN(n6) );
  LVT_IOA21HSV4 U2 ( .A1(n2), .A2(n4), .B(n5), .ZN(t_i_out) );
  LVT_INHSV2 U4 ( .I(n6), .ZN(n4) );
  LVT_INHSV2 U5 ( .I(n8), .ZN(n2) );
  LVT_NAND2HSV2 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U7 ( .A1(n8), .A2(n6), .ZN(n5) );
endmodule


module row_other_62 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_62 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_448 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_447 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_446 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_445 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_444 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_443 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_442 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_61 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_441 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_NAND2HSV2 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV1 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_440 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_439 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_438 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_CLKAND2HSV2 U1 ( .A1(b_in), .A2(a_in), .Z(n3) );
  LVT_XNOR2HSV4 U2 ( .A1(n3), .A2(t_i_1_in), .ZN(n4) );
  LVT_XOR2HSV2 U3 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_437 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_436 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_435 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U4 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV0P5 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2 U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_61 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_61 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_441 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_440 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_439 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_438 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_437 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_436 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_435 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_60 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_434 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_433 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_432 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_431 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_430 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .Z(n3) );
  LVT_XNOR2HSV4 U4 ( .A1(n3), .A2(t_i_1_in), .ZN(n4) );
endmodule


module cell_3_429 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_428 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV3SR U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV4 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV3SR U7 ( .I(n9), .ZN(n2) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_60 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_60 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_434 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_433 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_432 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_431 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_430 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_429 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_428 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_59 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_427 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_426 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_425 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_424 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_423 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_422 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKXOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_421 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV1 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV0 U4 ( .A1(n8), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U5 ( .I(t_i_1_in), .ZN(n4) );
  LVT_NAND2HSV2 U6 ( .A1(n5), .A2(n6), .ZN(n7) );
  LVT_INHSV2 U7 ( .I(n8), .ZN(n2) );
  LVT_XNOR2HSV4 U8 ( .A1(n9), .A2(n7), .ZN(t_i_out) );
endmodule


module row_other_59 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_59 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_427 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_426 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_425 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_424 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_423 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_422 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_421 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_58 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_420 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_419 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_418 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_417 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_416 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_415 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_414 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNHSV2 U2 ( .I(t_i_1_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(n8), .A2(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U6 ( .A1(n5), .A2(n6), .ZN(n7) );
  LVT_INHSV2 U7 ( .I(n8), .ZN(n2) );
  LVT_XNOR2HSV4 U8 ( .A1(n9), .A2(n7), .ZN(t_i_out) );
endmodule


module row_other_58 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_58 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_420 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_419 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_418 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_417 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_416 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_415 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_414 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_57 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n3), .A2(n4), .Z(t_i_out) );
endmodule


module cell_3_413 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_CLKXOR2HSV2 U1 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_XNOR2HSV1 U2 ( .A1(t_i_1_in), .A2(n3), .ZN(n4) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKAND2HSV2 U4 ( .A1(b_in), .A2(a_in), .Z(n3) );
endmodule


module cell_3_412 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_411 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_410 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_409 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_408 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_407 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(n8), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV2 U2 ( .I(t_i_1_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U5 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV2 U6 ( .A1(n5), .A2(n6), .ZN(n7) );
  LVT_INHSV2 U7 ( .I(n8), .ZN(n2) );
  LVT_XNOR2HSV4 U8 ( .A1(n9), .A2(n7), .ZN(t_i_out) );
endmodule


module row_other_57 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_57 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_413 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_412 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_411 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_410 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_409 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_408 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_407 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_56 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_406 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_405 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U5 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0P5 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_404 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_OAI21HSV2 U1 ( .A1(n6), .A2(n9), .B(n7), .ZN(t_i_out) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n9) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n9), .ZN(n7) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U6 ( .I(n8), .ZN(n4) );
  LVT_CLKNHSV2 U7 ( .I(n10), .ZN(n6) );
  LVT_NAND2HSV0P5 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_403 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_402 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10, n11;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n9) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n10) );
  LVT_INAND2HSV2 U2 ( .A1(n11), .B1(n10), .ZN(n8) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U5 ( .I(n9), .ZN(n4) );
  LVT_NAND2HSV0P5 U6 ( .A1(n11), .A2(n6), .ZN(n7) );
  LVT_NAND2HSV1 U7 ( .A1(n7), .A2(n8), .ZN(t_i_out) );
  LVT_INHSV0SR U8 ( .I(n10), .ZN(n6) );
  LVT_NAND2HSV0P5 U9 ( .A1(t_m_1_in), .A2(g_in), .ZN(n11) );
endmodule


module cell_3_401 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_400 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNHSV2 U4 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV0 U5 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV1 U6 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNHSV2 U7 ( .I(n9), .ZN(n2) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_56 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_56 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_406 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_405 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_404 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_403 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_402 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_401 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_400 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_8 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_8 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), .t_i_1_out(t0), 
        .t_i_2_out(t_i_2_out[6]) );
  row_other_62 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_61 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_60 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_59 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_58 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_57 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_56 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_49 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_48 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_7bit_32 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
endmodule


module PE_8 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   n22, l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1,
         n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n17, n18, n19, n20, n21
;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  LVT_NOR3HSV0 U24 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), .ZN(n18) );
  regist_8bit_53 u0 ( .clk(clk), .rstn(n15), .in(a_in), .out(l_a) );
  regist_8bit_52 u1 ( .clk(clk), .rstn(n15), .in(b_in), .out(b_out) );
  regist_8bit_51 u2 ( .clk(clk), .rstn(n15), .in(g_in), .out(l_g) );
  regist_1bit_35 u3 ( .clk(clk), .rstn(n15), .in(ctr), .out(l_ctr) );
  regist_1bit_34 u4 ( .clk(clk), .rstn(n15), .in(n11), .out(ctro) );
  regist_7bit_35 u5 ( .clk(clk), .rstn(n15), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_7bit_34 u6 ( .clk(clk), .rstn(n15), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_33 u7 ( .clk(clk), .rstn(n15), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_8bit_50 u9 ( .clk(clk), .rstn(n15), .in(mux_b), .out(mux_bq) );
  regist_1bit_32 u10 ( .clk(clk), .rstn(n15), .in(to_1), .out(ti_1) );
  regist_7bit_33 u11 ( .clk(clk), .rstn(n15), .in(to_7), .out(ti_7) );
  PE_core_8 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out({n22, t_i_2_out[5:0]}), .t_i_1_out_0(
        t_i_1_out_0) );
  regist_8bit_49 u12 ( .clk(clk), .rstn(n15), .in(ao), .out(a_out) );
  regist_8bit_48 u13 ( .clk(clk), .rstn(n15), .in(go), .out(g_out) );
  regist_7bit_32 u14 ( .clk(clk), .rstn(n15), .in(to), .out(t_i_1_out) );
  LVT_NOR4HSV4 U2 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(l_t_i_1_in[4]), 
        .A4(l_t_i_1_in[3]), .ZN(n17) );
  LVT_NAND2HSV2 U3 ( .A1(ti_7[0]), .A2(ctro), .ZN(n12) );
  LVT_CLKNAND2HSV4 U4 ( .A1(n7), .A2(n8), .ZN(to_7[2]) );
  LVT_NOR2HSV2 U5 ( .A1(n20), .A2(n19), .ZN(c_t_i_1_in_0) );
  LVT_NAND2HSV4 U6 ( .A1(t_i_2_out[0]), .A2(n21), .ZN(n13) );
  LVT_CLKNAND2HSV8 U7 ( .A1(n13), .A2(n12), .ZN(to_7[0]) );
  LVT_NAND2HSV4 U8 ( .A1(t_i_2_out[2]), .A2(n21), .ZN(n8) );
  LVT_AOI21HSV2 U9 ( .A1(n18), .A2(n17), .B(n6), .ZN(\c_t_i_1_in[0] ) );
  LVT_CLKNAND2HSV8 U10 ( .A1(n9), .A2(n10), .ZN(to_7[5]) );
  LVT_BUFHSV2 U11 ( .I(n19), .Z(n6) );
  LVT_INHSV0SR U12 ( .I(l_ctr), .ZN(n19) );
  LVT_INHSV2 U13 ( .I(ctro), .ZN(n21) );
  LVT_INHSV2 U14 ( .I(l_t_i_1_in_0), .ZN(n20) );
  LVT_AO22HSV2 U15 ( .A1(mux_bq[6]), .A2(l_ctr), .B1(b_out[6]), .B2(n6), .Z(
        mux_b[6]) );
  LVT_AO22HSV1 U16 ( .A1(mux_bq[1]), .A2(n11), .B1(b_out[1]), .B2(n6), .Z(
        mux_b[1]) );
  LVT_NAND2HSV2 U17 ( .A1(ti_7[2]), .A2(ctro), .ZN(n7) );
  LVT_NAND2HSV0P5 U18 ( .A1(ti_7[5]), .A2(ctro), .ZN(n9) );
  LVT_CLKNAND2HSV4 U19 ( .A1(t_i_2_out[5]), .A2(n21), .ZN(n10) );
  LVT_INHSV6 U20 ( .I(n16), .ZN(n15) );
  LVT_CLKNHSV1 U21 ( .I(n6), .ZN(n11) );
  LVT_AO22HSV2 U22 ( .A1(mux_bq[5]), .A2(l_ctr), .B1(b_out[5]), .B2(n6), .Z(
        mux_b[5]) );
  LVT_AO22HSV2 U23 ( .A1(mux_bq[4]), .A2(n11), .B1(b_out[4]), .B2(n6), .Z(
        mux_b[4]) );
  LVT_AO22HSV2 U25 ( .A1(mux_bq[3]), .A2(n11), .B1(b_out[3]), .B2(n6), .Z(
        mux_b[3]) );
  LVT_AO22HSV2 U26 ( .A1(mux_bq[7]), .A2(l_ctr), .B1(b_out[7]), .B2(n6), .Z(
        mux_b[7]) );
  LVT_AO22HSV2 U27 ( .A1(mux_bq[2]), .A2(n11), .B1(b_out[2]), .B2(n6), .Z(
        mux_b[2]) );
  LVT_AO22HSV2 U28 ( .A1(mux_bq[0]), .A2(n11), .B1(b_out[0]), .B2(n6), .Z(
        mux_b[0]) );
  LVT_BUFHSV2RT U29 ( .I(n22), .Z(t_i_2_out[6]) );
  LVT_AO22HSV4 U30 ( .A1(ti_7[1]), .A2(ctro), .B1(t_i_2_out[1]), .B2(n21), .Z(
        to_7[1]) );
  LVT_AO22HSV4 U31 ( .A1(ti_7[3]), .A2(ctro), .B1(t_i_2_out[3]), .B2(n21), .Z(
        to_7[3]) );
  LVT_AO22HSV4 U32 ( .A1(ti_7[4]), .A2(ctro), .B1(t_i_2_out[4]), .B2(n21), .Z(
        to_7[4]) );
  LVT_AO22HSV4 U33 ( .A1(ti_7[6]), .A2(ctro), .B1(n22), .B2(n21), .Z(to_7[6])
         );
  LVT_MOAI22HSV4 U34 ( .A1(l_ctr), .A2(n20), .B1(ti_1), .B2(l_ctr), .ZN(to_1)
         );
  LVT_INHSV2 U35 ( .I(rstn), .ZN(n16) );
endmodule


module regist_8bit_47 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_46 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_45 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_31 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_30 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV1 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_31 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV4 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV4 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV4 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_30 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
endmodule


module regist_1bit_29 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_44 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_28 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_29 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module cell_3_399 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_55 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_XOR2HSV2 U2 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKNAND2HSV1 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV2 U5 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_54 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_53 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U3 ( .A1(n5), .A2(n6), .Z(n7) );
endmodule


module cell_4_52 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n2), .A3(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_NAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_4_51 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV2 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_50 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_OAI21HSV2 U1 ( .A1(n5), .A2(n9), .B(n6), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n7) );
  LVT_XOR2HSV0 U3 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n10) );
  LVT_CLKXOR2HSV2 U5 ( .A1(n7), .A2(n8), .Z(n9) );
  LVT_NAND2HSV0P5 U6 ( .A1(n5), .A2(n9), .ZN(n6) );
  LVT_INHSV0SR U7 ( .I(n10), .ZN(n5) );
endmodule


module cell_4_49 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n2, n5, n6, n7, n8, n9, n10;

  LVT_INAND2HSV2 U1 ( .A1(n10), .B1(n9), .ZN(n6) );
  LVT_IOA21HSV2 U2 ( .A1(n6), .A2(n7), .B(n8), .ZN(n1) );
  LVT_INAND3HSV1 U3 ( .A1(n8), .B1(n6), .B2(n7), .ZN(n2) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U5 ( .A1(n5), .A2(n10), .ZN(n7) );
  LVT_NAND2HSV0P5 U6 ( .A1(b_in), .A2(a_in), .ZN(n10) );
  LVT_INHSV2 U7 ( .I(n9), .ZN(n5) );
  LVT_XNOR2HSV1 U8 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n8) );
  LVT_NAND2HSV2 U9 ( .A1(n1), .A2(n2), .ZN(t_i_out) );
endmodule


module row_1_7 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_3_399 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_55 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(t_i_1_out[1])
         );
  cell_4_54 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_53 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(
        t_i_1_out[3]) );
  cell_4_52 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(
        t_i_1_out[4]) );
  cell_4_51 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(
        t_i_1_out[5]) );
  cell_4_50 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_49 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
  LVT_CLKNHSV2 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_55 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_398 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_397 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_396 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U2 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_395 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_394 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_393 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_INAND2HSV2 U1 ( .A1(n8), .B1(n2), .ZN(n5) );
  LVT_CLKNHSV0 U2 ( .I(n6), .ZN(n2) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(n5), .ZN(t_i_out) );
  LVT_NAND2HSV0 U5 ( .A1(n6), .A2(n8), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XNOR2HSV4 U7 ( .A1(n7), .A2(t_i_1_in), .ZN(n6) );
endmodule


module cell_3_392 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U4 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV3 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2SR U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_55 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_55 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_398 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_397 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_396 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_395 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_394 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_393 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_392 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV1 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_54 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_391 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_390 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_389 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_388 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_XNOR2HSV1 U3 ( .A1(t_i_1_in), .A2(n3), .ZN(n4) );
  LVT_CLKAND2HSV2 U4 ( .A1(b_in), .A2(a_in), .Z(n3) );
endmodule


module cell_3_387 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_386 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_385 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV2 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U4 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV4 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV1 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2SR U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_54 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_54 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_391 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_390 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_389 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_388 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_387 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_386 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_385 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_53 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_384 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_383 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_382 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_381 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_NAND2HSV0 U1 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U3 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_380 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_379 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_378 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV2 U2 ( .A1(t_i_1_in), .A2(n8), .ZN(n5) );
  LVT_NAND2HSV2 U4 ( .A1(n5), .A2(n6), .ZN(n7) );
  LVT_INHSV2 U5 ( .I(t_i_1_in), .ZN(n2) );
  LVT_INHSV2 U6 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV4 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV4 U8 ( .A1(n9), .A2(n7), .ZN(t_i_out) );
endmodule


module row_other_53 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_53 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_384 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_383 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_382 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_381 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_380 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_379 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_378 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_52 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_377 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_376 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_375 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n12) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n14) );
  LVT_NAND2HSV2 U2 ( .A1(n12), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U5 ( .A1(n6), .A2(n7), .ZN(n13) );
  LVT_INHSV0SR U6 ( .I(n12), .ZN(n4) );
  LVT_INHSV2 U7 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV2 U8 ( .A1(n8), .A2(n13), .ZN(n11) );
  LVT_NAND2HSV0P5 U9 ( .A1(n14), .A2(n9), .ZN(n10) );
  LVT_NAND2HSV2 U10 ( .A1(n10), .A2(n11), .ZN(t_i_out) );
  LVT_INHSV0P5 U11 ( .I(n14), .ZN(n8) );
  LVT_INHSV2SR U12 ( .I(n13), .ZN(n9) );
endmodule


module cell_3_374 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_373 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_372 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_371 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U5 ( .I(n9), .ZN(n2) );
  LVT_INHSV2 U6 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV0 U7 ( .A1(n7), .A2(n9), .ZN(n5) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_52 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_52 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_377 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_376 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_375 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_374 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_373 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_372 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_371 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_51 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n3), .A2(n4), .Z(t_i_out) );
endmodule


module cell_3_370 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_369 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_368 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_367 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_NAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_366 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_365 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_364 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV2SR U2 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U5 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U6 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV0P5 U7 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_51 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_51 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_370 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_369 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_368 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_367 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_366 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_365 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_364 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_50 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_363 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_362 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_361 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_360 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_359 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_358 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_357 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module row_other_50 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_50 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_363 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_362 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_361 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_360 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_359 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_358 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_357 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_49 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4, n5, n6, n7;

  LVT_INAND2HSV2 U1 ( .A1(n6), .B1(n7), .ZN(n4) );
  LVT_NAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(n3), .A2(n6), .ZN(n5) );
  LVT_NAND2HSV0 U4 ( .A1(n4), .A2(n5), .ZN(t_i_out) );
  LVT_CLKNHSV0 U5 ( .I(n7), .ZN(n3) );
  LVT_NAND2HSV0P5 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_356 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_355 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_INAND2HSV2 U1 ( .A1(n9), .B1(n8), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n7), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKNAND2HSV0 U4 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV0P5 U6 ( .A1(n9), .A2(n4), .ZN(n5) );
  LVT_INHSV0SR U7 ( .I(n8), .ZN(n4) );
endmodule


module cell_3_354 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV2 U2 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U5 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV2 U6 ( .I(n8), .ZN(n4) );
  LVT_INHSV2 U7 ( .I(t_i_1_in), .ZN(n5) );
  LVT_CLKXOR2HSV2 U8 ( .A1(n10), .A2(n9), .Z(t_i_out) );
endmodule


module cell_3_353 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKXOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_352 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_351 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_350 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module row_other_49 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_49 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_356 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_355 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_354 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_353 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_352 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_351 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_350 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_7 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;
  wire   n1;
  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_7 u0 ( .a_in(a_in), .g_in({g_out[7], g_in[6:0]}), .b_in(b_in[7]), 
        .t_m_1_in(t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(
        t_i_2_in), .t_i_1_out(t0), .t_i_2_out(t_i_2_out[6]) );
  row_other_55 u1 ( .a_in(a_in), .g_in({g_out[7], g_in[6:0]}), .b_in(b_in[6]), 
        .t_m_1_in(t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(
        t_i_2_out[5]) );
  row_other_54 u2 ( .a_in(a_in), .g_in({g_out[7], g_in[6:0]}), .b_in(b_in[5]), 
        .t_m_1_in(t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(
        t_i_2_out[4]) );
  row_other_53 u3 ( .a_in(a_in), .g_in({g_out[7], g_in[6:0]}), .b_in(b_in[4]), 
        .t_m_1_in(t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(
        t_i_2_out[3]) );
  row_other_52 u4 ( .a_in(a_in), .g_in({g_out[7], g_in[6:0]}), .b_in(b_in[3]), 
        .t_m_1_in(t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(
        t_i_2_out[2]) );
  row_other_51 u5 ( .a_in(a_in), .g_in({g_out[7], g_in[6:0]}), .b_in(b_in[2]), 
        .t_m_1_in(t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(
        t_i_2_out[1]) );
  row_other_50 u6 ( .a_in(a_in), .g_in({g_out[7], g_in[6:0]}), .b_in(b_in[1]), 
        .t_m_1_in(t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(
        t_i_2_out[0]) );
  row_other_49 u7 ( .a_in(a_in), .g_in({g_out[7], g_in[6:0]}), .b_in(b_in[0]), 
        .t_m_1_in(t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), 
        .t_i_2_out(t_i_1_out_0) );
  LVT_INHSV2 U1 ( .I(g_in[7]), .ZN(n1) );
  LVT_INHSV4 U2 ( .I(n1), .ZN(g_out[7]) );
endmodule


module regist_8bit_43 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_42 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_7bit_28 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
endmodule


module PE_7 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  LVT_NOR3HSV0 U24 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), .ZN(n17) );
  regist_8bit_47 u0 ( .clk(clk), .rstn(n14), .in(a_in), .out(l_a) );
  regist_8bit_46 u1 ( .clk(clk), .rstn(n14), .in(b_in), .out(b_out) );
  regist_8bit_45 u2 ( .clk(clk), .rstn(n14), .in(g_in), .out(l_g) );
  regist_1bit_31 u3 ( .clk(clk), .rstn(n14), .in(ctr), .out(l_ctr) );
  regist_1bit_30 u4 ( .clk(clk), .rstn(n14), .in(n13), .out(ctro) );
  regist_7bit_31 u5 ( .clk(clk), .rstn(n14), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_7bit_30 u6 ( .clk(clk), .rstn(n14), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_29 u7 ( .clk(clk), .rstn(n14), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_8bit_44 u9 ( .clk(clk), .rstn(n14), .in(mux_b), .out(mux_bq) );
  regist_1bit_28 u10 ( .clk(clk), .rstn(n14), .in(to_1), .out(ti_1) );
  regist_7bit_29 u11 ( .clk(clk), .rstn(n14), .in(to_7), .out(ti_7) );
  PE_core_7 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out(t_i_2_out), .t_i_1_out_0(t_i_1_out_0)
         );
  regist_8bit_43 u12 ( .clk(clk), .rstn(n14), .in(ao), .out(a_out) );
  regist_8bit_42 u13 ( .clk(clk), .rstn(n14), .in(go), .out(g_out) );
  regist_7bit_28 u14 ( .clk(clk), .rstn(n14), .in(to), .out(t_i_1_out) );
  LVT_CLKNHSV4 U2 ( .I(l_t_i_1_in_0), .ZN(n19) );
  LVT_NOR3HSV12 U3 ( .A1(l_t_i_1_in[3]), .A2(l_t_i_1_in[5]), .A3(l_t_i_1_in[6]), .ZN(n7) );
  LVT_NOR2HSV2 U4 ( .A1(n19), .A2(n18), .ZN(c_t_i_1_in_0) );
  LVT_NAND2HSV4 U5 ( .A1(t_i_2_out[6]), .A2(n20), .ZN(n10) );
  LVT_INHSV3SR U6 ( .I(n7), .ZN(n8) );
  LVT_NAND2HSV8 U7 ( .A1(n12), .A2(n11), .ZN(to_7[2]) );
  LVT_BUFHSV2 U8 ( .I(n18), .Z(n6) );
  LVT_INHSV0SR U9 ( .I(l_ctr), .ZN(n18) );
  LVT_AOI21HSV0 U10 ( .A1(n17), .A2(n16), .B(n6), .ZN(\c_t_i_1_in[0] ) );
  LVT_NAND2HSV4 U11 ( .A1(t_i_2_out[2]), .A2(n20), .ZN(n12) );
  LVT_CLKNAND2HSV4 U12 ( .A1(n9), .A2(n10), .ZN(to_7[6]) );
  LVT_NAND2HSV2 U13 ( .A1(ti_7[2]), .A2(ctro), .ZN(n11) );
  LVT_AO22HSV1 U14 ( .A1(mux_bq[0]), .A2(n13), .B1(b_out[0]), .B2(n6), .Z(
        mux_b[0]) );
  LVT_AO22HSV1 U15 ( .A1(mux_bq[1]), .A2(n13), .B1(b_out[1]), .B2(n6), .Z(
        mux_b[1]) );
  LVT_AO22HSV1 U16 ( .A1(mux_bq[2]), .A2(n13), .B1(b_out[2]), .B2(n6), .Z(
        mux_b[2]) );
  LVT_AO22HSV1 U17 ( .A1(mux_bq[3]), .A2(n13), .B1(b_out[3]), .B2(n6), .Z(
        mux_b[3]) );
  LVT_AO22HSV1 U18 ( .A1(mux_bq[4]), .A2(n13), .B1(b_out[4]), .B2(n6), .Z(
        mux_b[4]) );
  LVT_AO22HSV1 U19 ( .A1(mux_bq[5]), .A2(n13), .B1(b_out[5]), .B2(n6), .Z(
        mux_b[5]) );
  LVT_AO22HSV1 U20 ( .A1(mux_bq[6]), .A2(n13), .B1(b_out[6]), .B2(n6), .Z(
        mux_b[6]) );
  LVT_AO22HSV1 U21 ( .A1(mux_bq[7]), .A2(n13), .B1(b_out[7]), .B2(n6), .Z(
        mux_b[7]) );
  LVT_NOR2HSV2 U22 ( .A1(l_t_i_1_in[4]), .A2(n8), .ZN(n16) );
  LVT_NAND2HSV2 U23 ( .A1(ti_7[6]), .A2(ctro), .ZN(n9) );
  LVT_INHSV2 U25 ( .I(ctro), .ZN(n20) );
  LVT_INHSV6 U26 ( .I(n15), .ZN(n14) );
  LVT_INHSV0SR U27 ( .I(n6), .ZN(n13) );
  LVT_AO22HSV4 U28 ( .A1(ti_7[0]), .A2(ctro), .B1(t_i_2_out[0]), .B2(n20), .Z(
        to_7[0]) );
  LVT_AO22HSV4 U29 ( .A1(ti_7[1]), .A2(ctro), .B1(t_i_2_out[1]), .B2(n20), .Z(
        to_7[1]) );
  LVT_AO22HSV4 U30 ( .A1(ti_7[3]), .A2(ctro), .B1(t_i_2_out[3]), .B2(n20), .Z(
        to_7[3]) );
  LVT_AO22HSV4 U31 ( .A1(ti_7[4]), .A2(ctro), .B1(t_i_2_out[4]), .B2(n20), .Z(
        to_7[4]) );
  LVT_AO22HSV4 U32 ( .A1(ti_7[5]), .A2(ctro), .B1(t_i_2_out[5]), .B2(n20), .Z(
        to_7[5]) );
  LVT_MOAI22HSV4 U33 ( .A1(l_ctr), .A2(n19), .B1(l_ctr), .B2(ti_1), .ZN(to_1)
         );
  LVT_INHSV2 U34 ( .I(rstn), .ZN(n15) );
endmodule


module regist_8bit_41 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_40 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_39 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_27 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_26 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_27 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV4 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV4 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV4 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_26 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
endmodule


module regist_1bit_25 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_38 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_24 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_25 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module cell_3_349 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_48 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_CLKNAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV2 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV4 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_47 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_XOR2HSV2 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_46 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV2 U1 ( .A1(n5), .A2(n2), .A3(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_45 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_XOR2HSV2 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_44 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n5, n6, n7;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n7), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U3 ( .A1(n5), .A2(n6), .ZN(n2) );
endmodule


module cell_4_43 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10;

  LVT_INAND2HSV0 U1 ( .A1(n9), .B1(n8), .ZN(n7) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U3 ( .A1(n6), .A2(n7), .ZN(n10) );
  LVT_INHSV2 U4 ( .I(n8), .ZN(n5) );
  LVT_XNOR2HSV4 U5 ( .A1(n10), .A2(n1), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U6 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n1) );
  LVT_NAND2HSV0P5 U7 ( .A1(n5), .A2(n9), .ZN(n6) );
  LVT_NAND2HSV0 U8 ( .A1(b_in), .A2(a_in), .ZN(n9) );
endmodule


module cell_4_42 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  LVT_NAND2HSV0 U1 ( .A1(n9), .A2(n13), .ZN(n10) );
  LVT_CLKNAND2HSV1 U2 ( .A1(n10), .A2(n11), .ZN(n15) );
  LVT_NAND2HSV2 U3 ( .A1(n8), .A2(n14), .ZN(n11) );
  LVT_INHSV2SR U4 ( .I(n15), .ZN(n1) );
  LVT_NAND2HSV2 U5 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_NAND2HSV2 U6 ( .A1(n1), .A2(n5), .ZN(n7) );
  LVT_CLKNAND2HSV2 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n13) );
  LVT_XNOR2HSV1 U8 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n12) );
  LVT_INHSV2 U9 ( .I(n13), .ZN(n8) );
  LVT_NAND2HSV2 U10 ( .A1(b_in), .A2(a_in), .ZN(n14) );
  LVT_CLKNAND2HSV0 U11 ( .A1(n15), .A2(n12), .ZN(n6) );
  LVT_INHSV2 U12 ( .I(n12), .ZN(n5) );
  LVT_INHSV0SR U13 ( .I(n14), .ZN(n9) );
endmodule


module row_1_6 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_3_349 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_48 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(
        t_i_1_out[1]) );
  cell_4_47 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_46 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(
        t_i_1_out[3]) );
  cell_4_45 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(
        t_i_1_out[4]) );
  cell_4_44 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(
        t_i_1_out[5]) );
  cell_4_43 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_42 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
endmodule


module cell_2_48 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_348 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_347 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_346 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_345 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_344 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_343 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_342 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV4SR U4 ( .I(n9), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV4 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV0P5 U7 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_48 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_48 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_348 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_347 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_346 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_345 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_344 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_343 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_342 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_47 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n3), .A2(n4), .Z(t_i_out) );
endmodule


module cell_3_341 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_340 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_339 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_338 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_337 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_336 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV0 U2 ( .A1(n8), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV1 U4 ( .I(t_i_1_in), .ZN(n4) );
  LVT_NAND2HSV2 U5 ( .A1(n5), .A2(n6), .ZN(n7) );
  LVT_INHSV2 U6 ( .I(n8), .ZN(n2) );
  LVT_NAND2HSV0 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV4 U8 ( .A1(n9), .A2(n7), .ZN(t_i_out) );
endmodule


module cell_3_335 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12;

  LVT_OAI21HSV2 U1 ( .A1(n8), .A2(t_i_1_in), .B(n9), .ZN(n11) );
  LVT_CLKNAND2HSV3 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n12) );
  LVT_INHSV2SR U3 ( .I(n12), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(n11), .ZN(n7) );
  LVT_CLKNAND2HSV1 U6 ( .A1(n8), .A2(t_i_1_in), .ZN(n9) );
  LVT_INHSV2SR U7 ( .I(n11), .ZN(n5) );
  LVT_CLKNAND2HSV1 U8 ( .A1(n12), .A2(n5), .ZN(n6) );
  LVT_INHSV2 U9 ( .I(n10), .ZN(n8) );
  LVT_NAND2HSV0 U10 ( .A1(b_in), .A2(a_in), .ZN(n10) );
endmodule


module row_other_47 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_47 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_341 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_340 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_339 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_338 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_337 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_336 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_335 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_46 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_334 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_333 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_332 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_331 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_330 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_NAND2HSV2 U1 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNHSV1 U2 ( .I(t_i_1_in), .ZN(n4) );
  LVT_NAND2HSV0 U3 ( .A1(n8), .A2(t_i_1_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n9), .A2(n7), .ZN(t_i_out) );
  LVT_NAND2HSV2 U5 ( .A1(n5), .A2(n6), .ZN(n7) );
  LVT_INHSV2 U6 ( .I(n8), .ZN(n2) );
  LVT_NAND2HSV2 U7 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
endmodule


module cell_3_329 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_328 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV2 U1 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV0 U2 ( .A1(n7), .A2(n9), .ZN(n5) );
  LVT_INHSV2 U4 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV4 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_46 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_46 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_334 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_333 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_332 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_331 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_330 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_329 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_328 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_45 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_327 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_326 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_325 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_324 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_323 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_322 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_321 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV2SR U1 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV2 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U5 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV2 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV0P5 U7 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_45 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_45 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_327 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_326 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_325 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_324 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_323 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_322 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_321 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_44 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_320 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_319 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_318 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_317 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_316 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_315 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_314 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV0 U4 ( .A1(n8), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV2 U5 ( .I(t_i_1_in), .ZN(n4) );
  LVT_NAND2HSV2 U6 ( .A1(n5), .A2(n6), .ZN(n7) );
  LVT_INHSV2 U7 ( .I(n8), .ZN(n2) );
  LVT_XNOR2HSV4 U8 ( .A1(n9), .A2(n7), .ZN(t_i_out) );
endmodule


module row_other_44 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_44 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_320 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_319 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_318 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_317 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_316 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_315 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_314 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_43 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_313 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_312 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_311 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_310 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_309 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_308 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_307 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV2 U5 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U6 ( .I(n9), .ZN(n2) );
  LVT_XNOR2HSV1 U7 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNHSV2 U8 ( .I(n7), .ZN(n4) );
endmodule


module row_other_43 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_43 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_313 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_312 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_311 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_310 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_309 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_308 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_307 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_42 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_306 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV1 U3 ( .A1(n3), .A2(t_i_1_in), .ZN(n4) );
  LVT_CLKAND2HSV2 U4 ( .A1(b_in), .A2(a_in), .Z(n3) );
endmodule


module cell_3_305 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_304 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_303 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_302 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_301 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_300 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module row_other_42 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_42 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_306 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_305 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_304 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_303 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_302 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_301 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_300 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_6 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_6 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), .t_i_1_out(t0), 
        .t_i_2_out(t_i_2_out[6]) );
  row_other_48 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_47 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_46 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_45 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_44 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_43 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_42 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_37 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_36 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_7bit_24 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module PE_6 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1, n3,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20
;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  LVT_AO22HSV0 U11 ( .A1(mux_bq[7]), .A2(n14), .B1(b_out[7]), .B2(n13), .Z(
        mux_b[7]) );
  LVT_AO22HSV0 U14 ( .A1(mux_bq[4]), .A2(n14), .B1(b_out[4]), .B2(n13), .Z(
        mux_b[4]) );
  LVT_AO22HSV0 U15 ( .A1(mux_bq[3]), .A2(n14), .B1(b_out[3]), .B2(n13), .Z(
        mux_b[3]) );
  LVT_AO22HSV0 U16 ( .A1(mux_bq[2]), .A2(n14), .B1(b_out[2]), .B2(n13), .Z(
        mux_b[2]) );
  LVT_AO22HSV0 U17 ( .A1(mux_bq[1]), .A2(n14), .B1(b_out[1]), .B2(n13), .Z(
        mux_b[1]) );
  LVT_AO22HSV0 U18 ( .A1(mux_bq[0]), .A2(n14), .B1(b_out[0]), .B2(n13), .Z(
        mux_b[0]) );
  regist_8bit_41 u0 ( .clk(clk), .rstn(n15), .in(a_in), .out(l_a) );
  regist_8bit_40 u1 ( .clk(clk), .rstn(n15), .in(b_in), .out(b_out) );
  regist_8bit_39 u2 ( .clk(clk), .rstn(n15), .in(g_in), .out(l_g) );
  regist_1bit_27 u3 ( .clk(clk), .rstn(n15), .in(ctr), .out(l_ctr) );
  regist_1bit_26 u4 ( .clk(clk), .rstn(n15), .in(n14), .out(ctro) );
  regist_7bit_27 u5 ( .clk(clk), .rstn(n15), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_7bit_26 u6 ( .clk(clk), .rstn(n15), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_25 u7 ( .clk(clk), .rstn(n15), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_8bit_38 u9 ( .clk(clk), .rstn(n15), .in(mux_b), .out(mux_bq) );
  regist_1bit_24 u10 ( .clk(clk), .rstn(n15), .in(to_1), .out(ti_1) );
  regist_7bit_25 u11 ( .clk(clk), .rstn(n15), .in(to_7), .out(ti_7) );
  PE_core_6 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out(t_i_2_out), .t_i_1_out_0(t_i_1_out_0)
         );
  regist_8bit_37 u12 ( .clk(clk), .rstn(n15), .in(ao), .out(a_out) );
  regist_8bit_36 u13 ( .clk(clk), .rstn(n15), .in(go), .out(g_out) );
  regist_7bit_24 u14 ( .clk(clk), .rstn(n15), .in(to), .out(t_i_1_out) );
  LVT_CLKNAND2HSV3 U2 ( .A1(t_i_2_out[0]), .A2(n20), .ZN(n8) );
  LVT_NAND2HSV8 U3 ( .A1(n10), .A2(n9), .ZN(to_7[2]) );
  LVT_CLKNAND2HSV3 U4 ( .A1(t_i_2_out[2]), .A2(n20), .ZN(n10) );
  LVT_CLKNAND2HSV3 U5 ( .A1(t_i_2_out[6]), .A2(n20), .ZN(n6) );
  LVT_INHSV4 U6 ( .I(l_t_i_1_in_0), .ZN(n19) );
  LVT_CLKNAND2HSV4 U7 ( .A1(n11), .A2(n12), .ZN(to_7[4]) );
  LVT_NAND2HSV2 U8 ( .A1(t_i_2_out[4]), .A2(n20), .ZN(n12) );
  LVT_INHSV2 U9 ( .I(ctro), .ZN(n20) );
  LVT_CLKNAND2HSV4 U10 ( .A1(n3), .A2(n6), .ZN(to_7[6]) );
  LVT_NAND2HSV2 U12 ( .A1(ti_7[6]), .A2(ctro), .ZN(n3) );
  LVT_NAND2HSV2 U13 ( .A1(ti_7[0]), .A2(ctro), .ZN(n7) );
  LVT_NAND2HSV4 U19 ( .A1(n8), .A2(n7), .ZN(to_7[0]) );
  LVT_CLKNAND2HSV1 U20 ( .A1(ti_7[2]), .A2(ctro), .ZN(n9) );
  LVT_NAND2HSV2 U21 ( .A1(ti_7[4]), .A2(ctro), .ZN(n11) );
  LVT_INHSV6 U22 ( .I(n16), .ZN(n15) );
  LVT_AOI21HSV2 U23 ( .A1(n18), .A2(n17), .B(n13), .ZN(\c_t_i_1_in[0] ) );
  LVT_INHSV2SR U24 ( .I(l_ctr), .ZN(n13) );
  LVT_NOR3HSV2 U25 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), .ZN(n18) );
  LVT_NOR2HSV2 U26 ( .A1(n19), .A2(n13), .ZN(c_t_i_1_in_0) );
  LVT_AO22HSV1 U27 ( .A1(mux_bq[5]), .A2(n14), .B1(b_out[5]), .B2(n13), .Z(
        mux_b[5]) );
  LVT_AO22HSV1 U28 ( .A1(mux_bq[6]), .A2(n14), .B1(b_out[6]), .B2(n13), .Z(
        mux_b[6]) );
  LVT_MOAI22HSV4 U29 ( .A1(l_ctr), .A2(n19), .B1(ti_1), .B2(l_ctr), .ZN(to_1)
         );
  LVT_NOR4HSV12 U30 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(
        l_t_i_1_in[4]), .A4(l_t_i_1_in[3]), .ZN(n17) );
  LVT_INHSV2 U31 ( .I(n13), .ZN(n14) );
  LVT_AO22HSV4 U32 ( .A1(ti_7[1]), .A2(ctro), .B1(t_i_2_out[1]), .B2(n20), .Z(
        to_7[1]) );
  LVT_AO22HSV4 U33 ( .A1(ti_7[3]), .A2(ctro), .B1(t_i_2_out[3]), .B2(n20), .Z(
        to_7[3]) );
  LVT_AO22HSV4 U34 ( .A1(ti_7[5]), .A2(ctro), .B1(t_i_2_out[5]), .B2(n20), .Z(
        to_7[5]) );
  LVT_INHSV2 U35 ( .I(rstn), .ZN(n16) );
endmodule


module regist_8bit_35 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_34 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_33 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_23 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_22 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV1 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_23 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_22 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
endmodule


module regist_1bit_21 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_32 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_20 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_21 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module cell_3_299 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_41 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_40 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U3 ( .A1(n7), .A2(n8), .Z(t_i_out) );
endmodule


module cell_4_39 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n2), .A3(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_38 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_37 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_36 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n9) );
  LVT_INAND2HSV2 U1 ( .A1(n10), .B1(n2), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n10) );
  LVT_INHSV2 U3 ( .I(n7), .ZN(n2) );
  LVT_XNOR2HSV1 U5 ( .A1(n8), .A2(n9), .ZN(n7) );
  LVT_NAND2HSV0P5 U6 ( .A1(n10), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV2 U7 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_4_35 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  LVT_INAND2HSV0 U1 ( .A1(n13), .B1(n12), .ZN(n10) );
  LVT_CLKNAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n12) );
  LVT_CLKNHSV2 U3 ( .I(n12), .ZN(n9) );
  LVT_NAND2HSV2 U4 ( .A1(n11), .A2(n10), .ZN(n14) );
  LVT_NAND2HSV2 U5 ( .A1(n9), .A2(n13), .ZN(n11) );
  LVT_INHSV2 U6 ( .I(n14), .ZN(n1) );
  LVT_CLKNAND2HSV1 U7 ( .A1(n8), .A2(n14), .ZN(n6) );
  LVT_NAND2HSV4 U8 ( .A1(n1), .A2(n5), .ZN(n7) );
  LVT_CLKNAND2HSV3 U9 ( .A1(n7), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV2 U10 ( .I(n8), .ZN(n5) );
  LVT_XNOR2HSV1 U11 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n8) );
  LVT_NAND2HSV0 U12 ( .A1(b_in), .A2(a_in), .ZN(n13) );
endmodule


module row_1_5 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_3_299 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_41 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(
        t_i_1_out[1]) );
  cell_4_40 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_39 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(
        t_i_1_out[3]) );
  cell_4_38 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(
        t_i_1_out[4]) );
  cell_4_37 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(
        t_i_1_out[5]) );
  cell_4_36 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_35 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_41 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_298 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_297 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_296 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_295 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_294 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_293 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  LVT_NAND2HSV2 U1 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .ZN(n12) );
  LVT_NAND2HSV0P5 U3 ( .A1(n14), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(n13), .ZN(n7) );
  LVT_INHSV2SR U5 ( .I(n14), .ZN(n4) );
  LVT_INHSV0SR U6 ( .I(n13), .ZN(n5) );
  LVT_NAND2HSV0P5 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n14) );
  LVT_NAND2HSV0P5 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n11) );
  LVT_CLKNHSV2 U9 ( .I(t_i_1_in), .ZN(n9) );
  LVT_NAND2HSV2 U10 ( .A1(n12), .A2(n9), .ZN(n10) );
  LVT_NAND2HSV2 U11 ( .A1(n10), .A2(n11), .ZN(n13) );
  LVT_CLKNHSV1 U12 ( .I(n12), .ZN(n8) );
endmodule


module cell_3_292 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV2 U2 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n7), .A2(n9), .ZN(n5) );
  LVT_INHSV4SR U6 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV4 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_41 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_41 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_298 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_297 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_296 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_295 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_294 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_293 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_292 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_40 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n3), .A2(n4), .Z(t_i_out) );
endmodule


module cell_3_291 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_290 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_289 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_288 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_287 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_286 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_285 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV3SR U1 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV0 U2 ( .A1(n7), .A2(n9), .ZN(n5) );
  LVT_CLKNHSV3 U4 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV4 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV4 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_40 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_40 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_291 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_290 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_289 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_288 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_287 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_286 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_285 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_39 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_284 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_283 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_CLKNHSV0P5 U6 ( .I(n8), .ZN(n4) );
endmodule


module cell_3_282 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_281 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_280 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_279 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_278 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV2SR U4 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV2 U5 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U6 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV0P5 U7 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2 U8 ( .I(n7), .ZN(n4) );
endmodule


module row_other_39 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_39 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_284 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_283 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_282 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_281 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_280 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_279 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_278 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_38 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n3), .A2(n4), .Z(t_i_out) );
endmodule


module cell_3_277 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_276 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_275 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_274 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_273 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_272 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKXOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_271 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV4SR U1 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV4 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_CLKNHSV4 U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV2 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV4 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_38 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_38 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_277 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_276 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_275 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_274 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_273 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_272 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_271 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_37 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_270 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_269 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_268 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_267 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_266 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_265 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_264 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV4SR U1 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV4 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV2 U4 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV0 U5 ( .A1(n7), .A2(n9), .ZN(n5) );
  LVT_NAND2HSV4 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U7 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
  LVT_CLKNAND2HSV3 U8 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
endmodule


module row_other_37 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_37 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_270 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_269 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_268 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_267 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_266 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_265 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_264 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_36 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_263 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_262 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_261 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_260 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_XNOR2HSV1 U3 ( .A1(t_i_1_in), .A2(n3), .ZN(n4) );
  LVT_CLKAND2HSV2 U4 ( .A1(b_in), .A2(a_in), .Z(n3) );
endmodule


module cell_3_259 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_258 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_257 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module row_other_36 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_36 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_263 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_262 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_261 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_260 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_259 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_258 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_257 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_35 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4, n5, n6, n7;

  LVT_INAND2HSV2 U1 ( .A1(n6), .B1(n7), .ZN(n4) );
  LVT_NAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_NAND2HSV1 U4 ( .A1(n4), .A2(n5), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U5 ( .A1(n3), .A2(n6), .ZN(n5) );
  LVT_INHSV2 U6 ( .I(n7), .ZN(n3) );
endmodule


module cell_3_256 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_XNOR2HSV1 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_255 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_INAND2HSV2 U1 ( .A1(n9), .B1(n8), .ZN(n6) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNHSV0P5 U4 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0P5 U5 ( .A1(n9), .A2(n4), .ZN(n5) );
  LVT_CLKNAND2HSV0 U6 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_XOR2HSV2 U7 ( .A1(n7), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_3_254 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_253 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV2 U1 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_CLKNHSV0P5 U2 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_CLKNAND2HSV0 U5 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_CLKNAND2HSV0 U6 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV0SR U7 ( .I(n10), .ZN(n4) );
  LVT_NAND2HSV0P5 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_252 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV1 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_251 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n8), .Z(n9) );
  LVT_INHSV0P5SR U2 ( .I(n10), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV0P5 U5 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U6 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_NAND2HSV0P5 U7 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_CLKNHSV1 U8 ( .I(n9), .ZN(n5) );
endmodule


module cell_3_250 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module row_other_35 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_35 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_256 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_255 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_254 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_253 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_252 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_251 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_250 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_5 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_5 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), .t_i_1_out(t0), 
        .t_i_2_out(t_i_2_out[6]) );
  row_other_41 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_40 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_39 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_38 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_37 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_36 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_35 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_31 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_30 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_7bit_20 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
endmodule


module PE_5 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  LVT_NOR3HSV0 U24 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), .ZN(n13) );
  regist_8bit_35 u0 ( .clk(clk), .rstn(n10), .in(a_in), .out(l_a) );
  regist_8bit_34 u1 ( .clk(clk), .rstn(n10), .in(b_in), .out(b_out) );
  regist_8bit_33 u2 ( .clk(clk), .rstn(n10), .in(g_in), .out(l_g) );
  regist_1bit_23 u3 ( .clk(clk), .rstn(n10), .in(ctr), .out(l_ctr) );
  regist_1bit_22 u4 ( .clk(clk), .rstn(n10), .in(n9), .out(ctro) );
  regist_7bit_23 u5 ( .clk(clk), .rstn(n10), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_7bit_22 u6 ( .clk(clk), .rstn(n10), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_21 u7 ( .clk(clk), .rstn(n10), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_8bit_32 u9 ( .clk(clk), .rstn(n10), .in(mux_b), .out(mux_bq) );
  regist_1bit_20 u10 ( .clk(clk), .rstn(n10), .in(n8), .out(ti_1) );
  regist_7bit_21 u11 ( .clk(clk), .rstn(n10), .in(to_7), .out(ti_7) );
  PE_core_5 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out(t_i_2_out), .t_i_1_out_0(t_i_1_out_0)
         );
  regist_8bit_31 u12 ( .clk(clk), .rstn(n10), .in(ao), .out(a_out) );
  regist_8bit_30 u13 ( .clk(clk), .rstn(n10), .in(go), .out(g_out) );
  regist_7bit_20 u14 ( .clk(clk), .rstn(n10), .in(to), .out(t_i_1_out) );
  LVT_INHSV0SR U2 ( .I(n14), .ZN(n9) );
  LVT_AO22HSV1 U3 ( .A1(mux_bq[4]), .A2(n9), .B1(b_out[4]), .B2(n14), .Z(
        mux_b[4]) );
  LVT_AO22HSV1 U4 ( .A1(mux_bq[3]), .A2(n9), .B1(b_out[3]), .B2(n14), .Z(
        mux_b[3]) );
  LVT_AO22HSV1 U5 ( .A1(mux_bq[2]), .A2(n9), .B1(b_out[2]), .B2(n14), .Z(
        mux_b[2]) );
  LVT_AO22HSV0 U6 ( .A1(mux_bq[7]), .A2(l_ctr), .B1(b_out[7]), .B2(n14), .Z(
        mux_b[7]) );
  LVT_AO22HSV0 U7 ( .A1(mux_bq[5]), .A2(l_ctr), .B1(b_out[5]), .B2(n14), .Z(
        mux_b[5]) );
  LVT_AO22HSV0 U8 ( .A1(mux_bq[6]), .A2(l_ctr), .B1(b_out[6]), .B2(n14), .Z(
        mux_b[6]) );
  LVT_CLKNAND2HSV4 U9 ( .A1(t_i_2_out[3]), .A2(n16), .ZN(n7) );
  LVT_CLKNAND2HSV8 U10 ( .A1(n7), .A2(n6), .ZN(to_7[3]) );
  LVT_AOI21HSV1 U11 ( .A1(n12), .A2(n13), .B(n14), .ZN(\c_t_i_1_in[0] ) );
  LVT_CLKNHSV1 U12 ( .I(l_ctr), .ZN(n14) );
  LVT_NOR4HSV12 U13 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(
        l_t_i_1_in[4]), .A4(l_t_i_1_in[3]), .ZN(n12) );
  LVT_AO22HSV1 U14 ( .A1(mux_bq[0]), .A2(n9), .B1(b_out[0]), .B2(n14), .Z(
        mux_b[0]) );
  LVT_AO22HSV1 U15 ( .A1(mux_bq[1]), .A2(n9), .B1(b_out[1]), .B2(n14), .Z(
        mux_b[1]) );
  LVT_NAND2HSV2 U16 ( .A1(ti_7[3]), .A2(ctro), .ZN(n6) );
  LVT_INHSV2 U17 ( .I(ctro), .ZN(n16) );
  LVT_INHSV4 U18 ( .I(l_t_i_1_in_0), .ZN(n15) );
  LVT_INHSV6 U19 ( .I(n11), .ZN(n10) );
  LVT_MOAI22HSV0 U20 ( .A1(l_ctr), .A2(n15), .B1(ti_1), .B2(l_ctr), .ZN(n8) );
  LVT_MOAI22HSV4 U21 ( .A1(l_ctr), .A2(n15), .B1(ti_1), .B2(l_ctr), .ZN(to_1)
         );
  LVT_NOR2HSV2 U22 ( .A1(n15), .A2(n14), .ZN(c_t_i_1_in_0) );
  LVT_AO22HSV4 U23 ( .A1(ti_7[0]), .A2(ctro), .B1(t_i_2_out[0]), .B2(n16), .Z(
        to_7[0]) );
  LVT_AO22HSV4 U25 ( .A1(ti_7[1]), .A2(ctro), .B1(t_i_2_out[1]), .B2(n16), .Z(
        to_7[1]) );
  LVT_AO22HSV4 U26 ( .A1(ti_7[2]), .A2(ctro), .B1(t_i_2_out[2]), .B2(n16), .Z(
        to_7[2]) );
  LVT_AO22HSV4 U27 ( .A1(ti_7[4]), .A2(ctro), .B1(t_i_2_out[4]), .B2(n16), .Z(
        to_7[4]) );
  LVT_AO22HSV4 U28 ( .A1(ti_7[5]), .A2(ctro), .B1(t_i_2_out[5]), .B2(n16), .Z(
        to_7[5]) );
  LVT_AO22HSV4 U29 ( .A1(ti_7[6]), .A2(ctro), .B1(t_i_2_out[6]), .B2(n16), .Z(
        to_7[6]) );
  LVT_INHSV2 U30 ( .I(rstn), .ZN(n11) );
endmodule


module regist_8bit_29 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_28 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_27 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_19 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_18 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_19 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV4 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV4 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_18 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_1bit_17 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_26 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_16 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_17 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module cell_3_249 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_34 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U3 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV2 U5 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_33 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_XOR2HSV2 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_32 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_31 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U3 ( .A1(n6), .A2(n5), .Z(n7) );
endmodule


module cell_4_30 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U3 ( .A1(n6), .A2(n5), .Z(n7) );
endmodule


module cell_4_29 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_XOR2HSV0 U1 ( .A1(n7), .A2(n6), .Z(n8) );
  LVT_OAI21HSV2 U2 ( .A1(n5), .A2(n8), .B(n1), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XNOR2HSV1 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U6 ( .A1(n5), .A2(n8), .ZN(n1) );
endmodule


module cell_4_28 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n13) );
  LVT_NAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .ZN(n14) );
  LVT_NAND2HSV1 U3 ( .A1(n15), .A2(n12), .ZN(n6) );
  LVT_CLKNAND2HSV0 U4 ( .A1(n9), .A2(n13), .ZN(n10) );
  LVT_NAND2HSV4 U5 ( .A1(n1), .A2(n5), .ZN(n7) );
  LVT_CLKNHSV2 U6 ( .I(n13), .ZN(n8) );
  LVT_XNOR2HSV1 U7 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n12) );
  LVT_CLKNAND2HSV3 U8 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV4SR U9 ( .I(n15), .ZN(n1) );
  LVT_INHSV2SR U10 ( .I(n12), .ZN(n5) );
  LVT_NAND2HSV4 U11 ( .A1(n10), .A2(n11), .ZN(n15) );
  LVT_CLKNAND2HSV3 U12 ( .A1(n8), .A2(n14), .ZN(n11) );
  LVT_INHSV0SR U13 ( .I(n14), .ZN(n9) );
endmodule


module row_1_4 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_3_249 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_34 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(
        t_i_1_out[1]) );
  cell_4_33 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_32 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(
        t_i_1_out[3]) );
  cell_4_31 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(
        t_i_1_out[4]) );
  cell_4_30 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(
        t_i_1_out[5]) );
  cell_4_29 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_28 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_34 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_248 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_247 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_246 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_245 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_244 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_243 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_242 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9, n10;

  LVT_OAI21HSV2 U1 ( .A1(t_i_1_in), .A2(n9), .B(n7), .ZN(n8) );
  LVT_CLKNAND2HSV2 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV0P5 U4 ( .A1(n10), .A2(n8), .ZN(n5) );
  LVT_NAND2HSV4 U5 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV3SR U6 ( .I(n10), .ZN(n2) );
  LVT_INHSV2 U7 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0P5 U8 ( .A1(n9), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV0 U9 ( .A1(b_in), .A2(a_in), .ZN(n9) );
endmodule


module row_other_34 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_34 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_248 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_247 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_246 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_245 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_244 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_243 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_242 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_33 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_241 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_240 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_239 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_238 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_237 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_236 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_CLKNHSV2 U2 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_XOR2HSV2 U5 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U6 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U7 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV2 U8 ( .I(n8), .ZN(n4) );
endmodule


module cell_3_235 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV4SR U2 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV1 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV4 U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV4 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_33 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_33 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_241 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_240 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_239 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_238 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_237 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_236 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_235 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_32 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_234 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_233 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_232 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_231 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_230 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_229 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_228 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U4 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV0 U5 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2 U6 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV2 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_32 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_32 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_234 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_233 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_232 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_231 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_230 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_229 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_228 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_31 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_227 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_226 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_225 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_224 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_223 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_222 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_221 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV2SR U1 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV0P5 U2 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV4 U5 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV2 U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_31 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_31 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_227 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_226 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_225 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_224 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_223 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_222 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_221 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_30 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n3), .A2(n4), .Z(t_i_out) );
endmodule


module cell_3_220 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_219 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_218 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_217 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_216 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_215 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_214 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module row_other_30 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_30 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_220 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_219 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_218 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_217 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_216 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_215 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_214 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_29 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n3), .A2(n4), .Z(t_i_out) );
endmodule


module cell_3_213 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_212 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_211 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_210 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_209 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_208 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_207 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV0 U2 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV3SR U4 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV4 U5 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV3SR U7 ( .I(n9), .ZN(n2) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_29 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_29 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_213 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_212 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_211 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_210 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_209 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_208 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_207 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_28 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n3), .A2(n4), .Z(t_i_out) );
endmodule


module cell_3_206 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_205 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_204 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n6), .Z(n7) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_INHSV1SR U5 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0P5 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_203 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_202 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_201 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_200 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKXOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module row_other_28 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_28 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_206 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_205 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_204 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_203 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_202 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_201 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_200 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_4 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_4 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), .t_i_1_out(t0), 
        .t_i_2_out(t_i_2_out[6]) );
  row_other_34 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_33 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_32 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_31 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_30 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_29 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_28 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_25 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_24 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_7bit_16 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
endmodule


module PE_4 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  regist_8bit_29 u0 ( .clk(clk), .rstn(n14), .in(a_in), .out(l_a) );
  regist_8bit_28 u1 ( .clk(clk), .rstn(n14), .in(b_in), .out(b_out) );
  regist_8bit_27 u2 ( .clk(clk), .rstn(n14), .in(g_in), .out(l_g) );
  regist_1bit_19 u3 ( .clk(clk), .rstn(n14), .in(ctr), .out(l_ctr) );
  regist_1bit_18 u4 ( .clk(clk), .rstn(n14), .in(n13), .out(ctro) );
  regist_7bit_19 u5 ( .clk(clk), .rstn(n14), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_7bit_18 u6 ( .clk(clk), .rstn(n14), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_17 u7 ( .clk(clk), .rstn(n14), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_8bit_26 u9 ( .clk(clk), .rstn(n14), .in(mux_b), .out(mux_bq) );
  regist_1bit_16 u10 ( .clk(clk), .rstn(n14), .in(n12), .out(ti_1) );
  regist_7bit_17 u11 ( .clk(clk), .rstn(n14), .in(to_7), .out(ti_7) );
  PE_core_4 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out(t_i_2_out), .t_i_1_out_0(t_i_1_out_0)
         );
  regist_8bit_25 u12 ( .clk(clk), .rstn(n14), .in(ao), .out(a_out) );
  regist_8bit_24 u13 ( .clk(clk), .rstn(n14), .in(go), .out(g_out) );
  regist_7bit_16 u14 ( .clk(clk), .rstn(n14), .in(to), .out(t_i_1_out) );
  LVT_AO22HSV1 U2 ( .A1(mux_bq[5]), .A2(n13), .B1(b_out[5]), .B2(n18), .Z(
        mux_b[5]) );
  LVT_AO22HSV1 U3 ( .A1(mux_bq[4]), .A2(n13), .B1(b_out[4]), .B2(n18), .Z(
        mux_b[4]) );
  LVT_AO22HSV1 U4 ( .A1(mux_bq[3]), .A2(n13), .B1(b_out[3]), .B2(n18), .Z(
        mux_b[3]) );
  LVT_AO22HSV1 U5 ( .A1(mux_bq[2]), .A2(n13), .B1(b_out[2]), .B2(n18), .Z(
        mux_b[2]) );
  LVT_AO22HSV1 U6 ( .A1(mux_bq[1]), .A2(n13), .B1(b_out[1]), .B2(n18), .Z(
        mux_b[1]) );
  LVT_INHSV2SR U7 ( .I(l_ctr), .ZN(n18) );
  LVT_INHSV3SR U8 ( .I(l_t_i_1_in_0), .ZN(n11) );
  LVT_INHSV2 U9 ( .I(ctro), .ZN(n20) );
  LVT_NAND2HSV2 U10 ( .A1(ti_7[4]), .A2(ctro), .ZN(n6) );
  LVT_CLKNAND2HSV4 U11 ( .A1(t_i_2_out[4]), .A2(n20), .ZN(n7) );
  LVT_NAND2HSV4 U12 ( .A1(n6), .A2(n7), .ZN(to_7[4]) );
  LVT_NAND2HSV0P5 U13 ( .A1(ti_7[2]), .A2(ctro), .ZN(n8) );
  LVT_CLKNAND2HSV4 U14 ( .A1(t_i_2_out[2]), .A2(n20), .ZN(n9) );
  LVT_NAND2HSV8 U15 ( .A1(n8), .A2(n9), .ZN(to_7[2]) );
  LVT_INHSV6 U16 ( .I(n15), .ZN(n14) );
  LVT_AOI21HSV2 U17 ( .A1(n17), .A2(n16), .B(n18), .ZN(\c_t_i_1_in[0] ) );
  LVT_NOR3HSV2 U18 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), .ZN(n17) );
  LVT_INHSV1SR U19 ( .I(n11), .ZN(n10) );
  LVT_INHSV0SR U20 ( .I(n10), .ZN(n19) );
  LVT_NOR2HSV1 U21 ( .A1(n19), .A2(n18), .ZN(c_t_i_1_in_0) );
  LVT_MOAI22HSV0 U22 ( .A1(n19), .A2(n13), .B1(ti_1), .B2(n13), .ZN(n12) );
  LVT_MOAI22HSV4 U23 ( .A1(n11), .A2(l_ctr), .B1(ti_1), .B2(l_ctr), .ZN(to_1)
         );
  LVT_INHSV0SR U24 ( .I(n18), .ZN(n13) );
  LVT_NOR4HSV12 U25 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(
        l_t_i_1_in[4]), .A4(l_t_i_1_in[3]), .ZN(n16) );
  LVT_AO22HSV2 U26 ( .A1(mux_bq[6]), .A2(n13), .B1(b_out[6]), .B2(n18), .Z(
        mux_b[6]) );
  LVT_AO22HSV2 U27 ( .A1(mux_bq[7]), .A2(n13), .B1(b_out[7]), .B2(n18), .Z(
        mux_b[7]) );
  LVT_AO22HSV2 U28 ( .A1(mux_bq[0]), .A2(n13), .B1(b_out[0]), .B2(n18), .Z(
        mux_b[0]) );
  LVT_AO22HSV4 U29 ( .A1(ti_7[0]), .A2(ctro), .B1(t_i_2_out[0]), .B2(n20), .Z(
        to_7[0]) );
  LVT_AO22HSV4 U30 ( .A1(ti_7[1]), .A2(ctro), .B1(t_i_2_out[1]), .B2(n20), .Z(
        to_7[1]) );
  LVT_AO22HSV4 U31 ( .A1(ti_7[3]), .A2(ctro), .B1(t_i_2_out[3]), .B2(n20), .Z(
        to_7[3]) );
  LVT_AO22HSV4 U32 ( .A1(ti_7[6]), .A2(ctro), .B1(t_i_2_out[6]), .B2(n20), .Z(
        to_7[6]) );
  LVT_AO22HSV4 U33 ( .A1(ti_7[5]), .A2(ctro), .B1(t_i_2_out[5]), .B2(n20), .Z(
        to_7[5]) );
  LVT_INHSV2 U34 ( .I(rstn), .ZN(n15) );
endmodule


module regist_8bit_23 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_22 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_21 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_15 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_14 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV1 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_15 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV4 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV4 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV4 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_14 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
endmodule


module regist_1bit_13 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_20 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_12 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_13 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module cell_3_199 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_27 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKXOR2HSV2 U3 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_XOR2HSV0 U5 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_26 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_XOR3HSV2 U2 ( .A1(n4), .A2(n2), .A3(n5), .Z(t_i_out) );
endmodule


module cell_4_25 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n5, n6, n7;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n7) );
  LVT_XNOR2HSV4 U1 ( .A1(n7), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n6), .ZN(n2) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_24 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_XOR3HSV1 U2 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
endmodule


module cell_4_23 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_XOR3HSV1 U2 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
endmodule


module cell_4_22 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8, n9, n10;

  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n10) );
  LVT_INAND2HSV2 U1 ( .A1(n7), .B1(n8), .ZN(n5) );
  LVT_INAND2HSV0 U2 ( .A1(n8), .B1(n7), .ZN(n6) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n7) );
  LVT_XOR2HSV4 U4 ( .A1(n9), .A2(n10), .Z(t_i_out) );
  LVT_NAND2HSV2 U6 ( .A1(n5), .A2(n6), .ZN(n9) );
  LVT_NAND2HSV0 U7 ( .A1(b_in), .A2(a_in), .ZN(n8) );
endmodule


module cell_4_21 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n13) );
  LVT_CLKNAND2HSV2 U2 ( .A1(n10), .A2(n14), .ZN(n11) );
  LVT_XNOR2HSV1 U3 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n8) );
  LVT_NAND2HSV1 U4 ( .A1(n8), .A2(n15), .ZN(n6) );
  LVT_CLKNAND2HSV3 U5 ( .A1(n11), .A2(n12), .ZN(n15) );
  LVT_NAND2HSV4 U6 ( .A1(n1), .A2(n5), .ZN(n7) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV3SR U8 ( .I(n15), .ZN(n1) );
  LVT_INHSV2SR U9 ( .I(n8), .ZN(n5) );
  LVT_CLKNHSV0P5 U10 ( .I(n13), .ZN(n10) );
  LVT_NAND2HSV0P5 U11 ( .A1(n9), .A2(n13), .ZN(n12) );
  LVT_INHSV0SR U12 ( .I(n14), .ZN(n9) );
  LVT_NAND2HSV0 U13 ( .A1(b_in), .A2(a_in), .ZN(n14) );
endmodule


module row_1_3 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_3_199 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_27 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(
        t_i_1_out[1]) );
  cell_4_26 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_25 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(
        t_i_1_out[3]) );
  cell_4_24 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(t_i_1_out[4])
         );
  cell_4_23 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(t_i_1_out[5])
         );
  cell_4_22 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_21 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
  LVT_INHSV2 U3 ( .I(n1), .ZN(n3) );
endmodule


module cell_2_27 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_198 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_197 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_196 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_195 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_194 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_193 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_192 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4, n5, n6, n7, n8;

  LVT_CLKXOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n6), .Z(n7) );
  LVT_CLKAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .Z(n6) );
  LVT_INHSV2 U3 ( .I(n7), .ZN(n3) );
  LVT_NAND2HSV4 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U5 ( .A1(n7), .A2(n8), .ZN(n4) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n4), .A2(n5), .ZN(t_i_out) );
  LVT_INHSV3SR U7 ( .I(n8), .ZN(n2) );
  LVT_NAND2HSV4 U8 ( .A1(n2), .A2(n3), .ZN(n5) );
endmodule


module row_other_27 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_27 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_198 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_197 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_196 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_195 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_194 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_193 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_192 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_26 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_191 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_190 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_189 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_188 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_187 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_186 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKXOR2HSV2 U1 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV4 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV0 U3 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNHSV0P5 U4 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV0P5 U5 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U6 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV2 U7 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV2 U8 ( .A1(b_in), .A2(a_in), .ZN(n8) );
endmodule


module cell_3_185 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module row_other_26 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_26 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_191 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_190 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_189 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_188 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_187 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_186 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_185 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_25 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_184 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_183 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_182 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_181 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_180 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_179 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_178 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4;

  LVT_CLKAND2HSV2 U1 ( .A1(b_in), .A2(a_in), .Z(n2) );
  LVT_XOR2HSV4 U2 ( .A1(t_i_1_in), .A2(n2), .Z(n3) );
  LVT_XNOR2HSV4 U3 ( .A1(n4), .A2(n3), .ZN(t_i_out) );
  LVT_NAND2HSV4 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n4) );
endmodule


module row_other_25 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_25 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_184 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_183 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_182 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_181 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_180 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_179 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_178 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_24 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_177 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_176 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_175 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_174 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_173 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_172 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_171 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_NAND2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNHSV0P5 U2 ( .I(t_i_1_in), .ZN(n5) );
  LVT_CLKXOR2HSV2 U3 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_NAND2HSV4 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV0P5 U6 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_INHSV2 U7 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0 U8 ( .A1(b_in), .A2(a_in), .ZN(n8) );
endmodule


module row_other_24 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_24 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_177 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_176 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_175 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_174 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_173 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_172 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_171 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_23 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(g_in), .A2(t_m_1_in), .ZN(n3) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_170 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_169 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_168 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_167 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_166 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_165 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_164 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XNOR2HSV1 U1 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
  LVT_INHSV2 U2 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV0P5 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNHSV4 U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV2 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV4 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U8 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
endmodule


module row_other_23 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_23 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_170 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_169 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_168 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_167 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_166 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_165 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_164 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_22 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_163 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV1 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_162 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_161 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_160 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_159 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_158 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_157 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(n7), .A2(n9), .ZN(n5) );
  LVT_INHSV4 U2 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
  LVT_INHSV3SR U5 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV2 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV4 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U8 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
endmodule


module row_other_22 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_22 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_163 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_162 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_161 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_160 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_159 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_158 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_157 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_21 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_156 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV1 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_155 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_154 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_153 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_152 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_151 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_150 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module row_other_21 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_21 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_156 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_155 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_154 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_153 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_152 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_151 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_150 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_3 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_3 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), .t_i_1_out(t0), 
        .t_i_2_out(t_i_2_out[6]) );
  row_other_27 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_26 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_25 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_24 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_23 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_22 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_21 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_19 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_18 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_7bit_12 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
endmodule


module PE_3 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  LVT_AO22HSV0 U13 ( .A1(mux_bq[5]), .A2(n10), .B1(b_out[5]), .B2(n17), .Z(
        mux_b[5]) );
  LVT_AO22HSV0 U14 ( .A1(mux_bq[4]), .A2(n10), .B1(b_out[4]), .B2(n17), .Z(
        mux_b[4]) );
  LVT_AO22HSV0 U15 ( .A1(mux_bq[3]), .A2(n10), .B1(b_out[3]), .B2(n17), .Z(
        mux_b[3]) );
  LVT_AO22HSV0 U16 ( .A1(mux_bq[2]), .A2(n10), .B1(b_out[2]), .B2(n17), .Z(
        mux_b[2]) );
  LVT_AO22HSV0 U17 ( .A1(mux_bq[1]), .A2(n10), .B1(b_out[1]), .B2(n17), .Z(
        mux_b[1]) );
  LVT_AO22HSV0 U18 ( .A1(mux_bq[0]), .A2(n10), .B1(b_out[0]), .B2(n17), .Z(
        mux_b[0]) );
  LVT_NOR2HSV0 U19 ( .A1(n18), .A2(n17), .ZN(c_t_i_1_in_0) );
  regist_8bit_23 u0 ( .clk(clk), .rstn(n13), .in(a_in), .out(l_a) );
  regist_8bit_22 u1 ( .clk(clk), .rstn(n13), .in(b_in), .out(b_out) );
  regist_8bit_21 u2 ( .clk(clk), .rstn(n13), .in(g_in), .out(l_g) );
  regist_1bit_15 u3 ( .clk(clk), .rstn(n13), .in(ctr), .out(l_ctr) );
  regist_1bit_14 u4 ( .clk(clk), .rstn(n13), .in(n10), .out(ctro) );
  regist_7bit_15 u5 ( .clk(clk), .rstn(n13), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_7bit_14 u6 ( .clk(clk), .rstn(n13), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_13 u7 ( .clk(clk), .rstn(n13), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_8bit_20 u9 ( .clk(clk), .rstn(n13), .in(mux_b), .out(mux_bq) );
  regist_1bit_12 u10 ( .clk(clk), .rstn(n13), .in(n9), .out(ti_1) );
  regist_7bit_13 u11 ( .clk(clk), .rstn(n13), .in(to_7), .out(ti_7) );
  PE_core_3 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out(t_i_2_out), .t_i_1_out_0(t_i_1_out_0)
         );
  regist_8bit_19 u12 ( .clk(clk), .rstn(n13), .in(ao), .out(a_out) );
  regist_8bit_18 u13 ( .clk(clk), .rstn(n13), .in(go), .out(g_out) );
  regist_7bit_12 u14 ( .clk(clk), .rstn(n13), .in(to), .out(t_i_1_out) );
  LVT_INHSV3SR U2 ( .I(l_t_i_1_in_0), .ZN(n18) );
  LVT_NAND2HSV2 U3 ( .A1(ti_7[4]), .A2(ctro), .ZN(n11) );
  LVT_INHSV2SR U4 ( .I(l_ctr), .ZN(n17) );
  LVT_CLKNAND2HSV4 U5 ( .A1(t_i_2_out[1]), .A2(n19), .ZN(n7) );
  LVT_NAND2HSV4 U6 ( .A1(t_i_2_out[4]), .A2(n19), .ZN(n12) );
  LVT_CLKNAND2HSV1 U7 ( .A1(ti_7[1]), .A2(ctro), .ZN(n6) );
  LVT_NAND2HSV8 U8 ( .A1(n7), .A2(n6), .ZN(to_7[1]) );
  LVT_INHSV2 U9 ( .I(ctro), .ZN(n19) );
  LVT_INHSV6 U10 ( .I(n14), .ZN(n13) );
  LVT_NOR3HSV2 U11 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), .ZN(n16) );
  LVT_NOR4HSV12 U12 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(
        l_t_i_1_in[4]), .A4(l_t_i_1_in[3]), .ZN(n15) );
  LVT_INHSV0SR U20 ( .I(to_1), .ZN(n8) );
  LVT_INHSV2 U21 ( .I(n8), .ZN(n9) );
  LVT_CLKNAND2HSV8 U22 ( .A1(n12), .A2(n11), .ZN(to_7[4]) );
  LVT_INHSV0SR U23 ( .I(n17), .ZN(n10) );
  LVT_AOI21HSV2 U24 ( .A1(n16), .A2(n15), .B(n17), .ZN(\c_t_i_1_in[0] ) );
  LVT_AO22HSV1 U25 ( .A1(mux_bq[6]), .A2(n10), .B1(b_out[6]), .B2(n17), .Z(
        mux_b[6]) );
  LVT_AO22HSV1 U26 ( .A1(mux_bq[7]), .A2(n10), .B1(b_out[7]), .B2(n17), .Z(
        mux_b[7]) );
  LVT_MOAI22HSV4 U27 ( .A1(n18), .A2(l_ctr), .B1(ti_1), .B2(l_ctr), .ZN(to_1)
         );
  LVT_AO22HSV4 U28 ( .A1(ti_7[0]), .A2(ctro), .B1(t_i_2_out[0]), .B2(n19), .Z(
        to_7[0]) );
  LVT_AO22HSV4 U29 ( .A1(ti_7[2]), .A2(ctro), .B1(t_i_2_out[2]), .B2(n19), .Z(
        to_7[2]) );
  LVT_AO22HSV4 U30 ( .A1(ti_7[3]), .A2(ctro), .B1(t_i_2_out[3]), .B2(n19), .Z(
        to_7[3]) );
  LVT_AO22HSV4 U31 ( .A1(ti_7[5]), .A2(ctro), .B1(t_i_2_out[5]), .B2(n19), .Z(
        to_7[5]) );
  LVT_AO22HSV4 U32 ( .A1(ti_7[6]), .A2(ctro), .B1(t_i_2_out[6]), .B2(n19), .Z(
        to_7[6]) );
  LVT_INHSV2 U33 ( .I(rstn), .ZN(n14) );
endmodule


module regist_8bit_17 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_16 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_15 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_11 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_10 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV1 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_11 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV4 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV4 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_10 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
endmodule


module regist_1bit_9 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_14 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_8 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_9 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module cell_3_149 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_20 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_XOR2HSV2 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_19 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(g_in), .A2(t_m_1_in), .ZN(n5) );
endmodule


module cell_4_18 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n2), .A3(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_17 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U1 ( .A1(g_in), .A2(t_m_1_in), .ZN(n2) );
  LVT_XOR3HSV1 U2 ( .A1(n5), .A2(n2), .A3(n4), .Z(t_i_out) );
endmodule


module cell_4_16 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n2), .A3(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_15 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n3, n4;

  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR3HSV1 U2 ( .A1(n4), .A2(n2), .A3(n3), .Z(t_i_out) );
  LVT_NAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .ZN(n2) );
endmodule


module cell_4_14 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  LVT_INHSV2 U1 ( .I(n13), .ZN(n10) );
  LVT_NAND2HSV0 U2 ( .A1(n9), .A2(n13), .ZN(n12) );
  LVT_CLKNAND2HSV1 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n13) );
  LVT_NAND2HSV2 U4 ( .A1(n11), .A2(n12), .ZN(n15) );
  LVT_NAND2HSV0P5 U5 ( .A1(n15), .A2(n8), .ZN(n6) );
  LVT_XNOR2HSV1 U6 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n8) );
  LVT_INHSV2 U7 ( .I(n15), .ZN(n1) );
  LVT_NAND2HSV0P5 U8 ( .A1(n10), .A2(n14), .ZN(n11) );
  LVT_CLKNAND2HSV3 U9 ( .A1(n1), .A2(n5), .ZN(n7) );
  LVT_CLKNAND2HSV3 U10 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV3SR U11 ( .I(n8), .ZN(n5) );
  LVT_INHSV0SR U12 ( .I(n14), .ZN(n9) );
  LVT_NAND2HSV0 U13 ( .A1(b_in), .A2(a_in), .ZN(n14) );
endmodule


module row_1_2 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_3_149 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_20 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(t_i_1_out[1])
         );
  cell_4_19 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_18 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(
        t_i_1_out[3]) );
  cell_4_17 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(
        t_i_1_out[4]) );
  cell_4_16 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(
        t_i_1_out[5]) );
  cell_4_15 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_14 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV0P5SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_20 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_148 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_147 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_146 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_145 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_144 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_143 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4;

  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n4) );
  LVT_CLKAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .Z(n2) );
  LVT_XOR2HSV0 U3 ( .A1(n2), .A2(t_i_1_in), .Z(n3) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(n3), .ZN(t_i_out) );
endmodule


module cell_3_142 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_XNOR2HSV1 U1 ( .A1(t_i_1_in), .A2(n7), .ZN(n6) );
  LVT_IOA21HSV4 U2 ( .A1(n2), .A2(n4), .B(n5), .ZN(t_i_out) );
  LVT_INHSV2 U4 ( .I(n6), .ZN(n4) );
  LVT_INHSV2 U5 ( .I(n8), .ZN(n2) );
  LVT_NAND2HSV2 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U7 ( .A1(n6), .A2(n8), .ZN(n5) );
endmodule


module row_other_20 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_20 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_148 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_147 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_146 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_145 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_144 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_143 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_142 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_19 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n3), .A2(n4), .Z(t_i_out) );
endmodule


module cell_3_141 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_140 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_139 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_138 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_CLKAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .Z(n3) );
  LVT_XNOR2HSV4 U4 ( .A1(n3), .A2(t_i_1_in), .ZN(n4) );
endmodule


module cell_3_137 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_136 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_135 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_NAND2HSV4 U1 ( .A1(n6), .A2(n4), .ZN(n2) );
  LVT_OAI21HSV2 U2 ( .A1(n6), .A2(n4), .B(n2), .ZN(t_i_out) );
  LVT_NAND2HSV4 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XNOR2HSV4 U5 ( .A1(n5), .A2(t_i_1_in), .ZN(n4) );
endmodule


module row_other_19 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_19 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_141 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_140 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_139 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_138 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_137 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_136 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_135 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_18 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_134 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_133 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_132 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_131 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_130 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_129 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_128 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0 U1 ( .A1(n8), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV0P5 U2 ( .I(t_i_1_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U6 ( .A1(n5), .A2(n6), .ZN(n7) );
  LVT_INHSV2 U7 ( .I(n8), .ZN(n2) );
  LVT_XNOR2HSV4 U8 ( .A1(n9), .A2(n7), .ZN(t_i_out) );
endmodule


module row_other_18 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_18 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_134 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_133 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_132 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_131 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_130 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_129 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_128 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_17 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_127 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_126 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_125 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_124 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_123 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_122 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5, n6;

  LVT_NAND2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n3) );
  LVT_OAI21HSV2 U2 ( .A1(t_i_1_in), .A2(n4), .B(n3), .ZN(n5) );
  LVT_NAND2HSV2 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKAND2HSV2 U4 ( .A1(b_in), .A2(a_in), .Z(n4) );
  LVT_XOR2HSV2 U5 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_121 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  LVT_NAND2HSV4 U1 ( .A1(n10), .A2(n11), .ZN(n13) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n12), .A2(n9), .ZN(n10) );
  LVT_INHSV2 U3 ( .I(n14), .ZN(n4) );
  LVT_NAND2HSV4 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n14) );
  LVT_CLKNAND2HSV3 U5 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_NAND2HSV2 U6 ( .A1(b_in), .A2(a_in), .ZN(n12) );
  LVT_INHSV3SR U7 ( .I(n13), .ZN(n5) );
  LVT_CLKNAND2HSV3 U8 ( .A1(n4), .A2(n13), .ZN(n7) );
  LVT_CLKNAND2HSV1 U9 ( .A1(n8), .A2(t_i_1_in), .ZN(n11) );
  LVT_CLKNHSV2P5 U10 ( .I(t_i_1_in), .ZN(n9) );
  LVT_NAND2HSV0P5 U11 ( .A1(n14), .A2(n5), .ZN(n6) );
  LVT_INHSV2 U12 ( .I(n12), .ZN(n8) );
endmodule


module row_other_17 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_17 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_127 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_126 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_125 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_124 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_123 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_122 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_121 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_16 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_120 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_119 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_118 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_117 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_116 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_115 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4;

  LVT_CLKXOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n3), .Z(n2) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(n2), .ZN(t_i_out) );
  LVT_CLKAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .Z(n3) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n4) );
endmodule


module cell_3_114 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV2SR U1 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV4 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n7), .A2(n9), .ZN(n5) );
  LVT_NAND2HSV4 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV4SR U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_16 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_16 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_120 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_119 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_118 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_117 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_116 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_115 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_114 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_15 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_113 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_112 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_111 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_110 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_109 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_108 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_107 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module row_other_15 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_15 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_113 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_112 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_111 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_110 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_109 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_108 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_107 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_14 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_106 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNHSV0P5 U1 ( .I(n10), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_NAND2HSV0P5 U4 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_CLKNAND2HSV0 U5 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_CLKNAND2HSV0 U6 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV0SR U7 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV0 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_105 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_104 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_103 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_102 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_101 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_100 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module row_other_14 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_14 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_106 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_105 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_104 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_103 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_102 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_101 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_100 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_2 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_2 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), .t_i_1_out(t0), 
        .t_i_2_out(t_i_2_out[6]) );
  row_other_20 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_19 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_18 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_17 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_16 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_15 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_14 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_13 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_12 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_7bit_8 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
endmodule


module PE_2 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  LVT_AOI21HSV0 U21 ( .A1(n17), .A2(n16), .B(n18), .ZN(\c_t_i_1_in[0] ) );
  LVT_NOR3HSV0 U24 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), .ZN(n17) );
  regist_8bit_17 u0 ( .clk(clk), .rstn(n14), .in(a_in), .out(l_a) );
  regist_8bit_16 u1 ( .clk(clk), .rstn(n14), .in(b_in), .out(b_out) );
  regist_8bit_15 u2 ( .clk(clk), .rstn(n14), .in(g_in), .out(l_g) );
  regist_1bit_11 u3 ( .clk(clk), .rstn(n14), .in(ctr), .out(l_ctr) );
  regist_1bit_10 u4 ( .clk(clk), .rstn(n14), .in(n11), .out(ctro) );
  regist_7bit_11 u5 ( .clk(clk), .rstn(n14), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_7bit_10 u6 ( .clk(clk), .rstn(n14), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_9 u7 ( .clk(clk), .rstn(n14), .in(t_i_1_in_0), .out(l_t_i_1_in_0) );
  regist_8bit_14 u9 ( .clk(clk), .rstn(n14), .in(mux_b), .out(mux_bq) );
  regist_1bit_8 u10 ( .clk(clk), .rstn(n14), .in(n10), .out(ti_1) );
  regist_7bit_9 u11 ( .clk(clk), .rstn(n14), .in(to_7), .out(ti_7) );
  PE_core_2 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out(t_i_2_out), .t_i_1_out_0(t_i_1_out_0)
         );
  regist_8bit_13 u12 ( .clk(clk), .rstn(n14), .in(ao), .out(a_out) );
  regist_8bit_12 u13 ( .clk(clk), .rstn(n14), .in(go), .out(g_out) );
  regist_7bit_8 u14 ( .clk(clk), .rstn(n14), .in(to), .out(t_i_1_out) );
  LVT_INHSV2 U2 ( .I(ctro), .ZN(n20) );
  LVT_INHSV1SR U3 ( .I(l_ctr), .ZN(n18) );
  LVT_NOR4HSV4 U4 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(l_t_i_1_in[4]), 
        .A4(l_t_i_1_in[3]), .ZN(n16) );
  LVT_NAND2HSV2 U5 ( .A1(ti_7[5]), .A2(ctro), .ZN(n6) );
  LVT_CLKNAND2HSV3 U6 ( .A1(t_i_2_out[5]), .A2(n20), .ZN(n7) );
  LVT_NAND2HSV4 U7 ( .A1(n6), .A2(n7), .ZN(to_7[5]) );
  LVT_NAND2HSV2 U8 ( .A1(ti_7[1]), .A2(ctro), .ZN(n8) );
  LVT_CLKNAND2HSV3 U9 ( .A1(t_i_2_out[1]), .A2(n20), .ZN(n9) );
  LVT_NAND2HSV4 U10 ( .A1(n8), .A2(n9), .ZN(to_7[1]) );
  LVT_INHSV6 U11 ( .I(n15), .ZN(n14) );
  LVT_IOA22HSV0 U12 ( .B1(l_ctr), .B2(n19), .A1(ti_1), .A2(l_ctr), .ZN(n10) );
  LVT_INHSV4 U13 ( .I(l_t_i_1_in_0), .ZN(n19) );
  LVT_MOAI22HSV4 U14 ( .A1(l_ctr), .A2(n19), .B1(ti_1), .B2(l_ctr), .ZN(to_1)
         );
  LVT_NOR2HSV0 U15 ( .A1(n19), .A2(n18), .ZN(c_t_i_1_in_0) );
  LVT_INHSV0SR U16 ( .I(n18), .ZN(n11) );
  LVT_CLKNAND2HSV8 U17 ( .A1(n12), .A2(n13), .ZN(to_7[3]) );
  LVT_NAND2HSV8 U18 ( .A1(t_i_2_out[3]), .A2(n20), .ZN(n13) );
  LVT_NAND2HSV4 U19 ( .A1(ti_7[3]), .A2(ctro), .ZN(n12) );
  LVT_AO22HSV2 U20 ( .A1(mux_bq[5]), .A2(n11), .B1(b_out[5]), .B2(n18), .Z(
        mux_b[5]) );
  LVT_AO22HSV2 U22 ( .A1(mux_bq[6]), .A2(n11), .B1(b_out[6]), .B2(n18), .Z(
        mux_b[6]) );
  LVT_AO22HSV2 U23 ( .A1(mux_bq[4]), .A2(n11), .B1(b_out[4]), .B2(n18), .Z(
        mux_b[4]) );
  LVT_AO22HSV2 U25 ( .A1(mux_bq[3]), .A2(n11), .B1(b_out[3]), .B2(n18), .Z(
        mux_b[3]) );
  LVT_AO22HSV2 U26 ( .A1(mux_bq[2]), .A2(n11), .B1(b_out[2]), .B2(n18), .Z(
        mux_b[2]) );
  LVT_AO22HSV2 U27 ( .A1(mux_bq[1]), .A2(n11), .B1(b_out[1]), .B2(n18), .Z(
        mux_b[1]) );
  LVT_AO22HSV2 U28 ( .A1(mux_bq[0]), .A2(n11), .B1(b_out[0]), .B2(n18), .Z(
        mux_b[0]) );
  LVT_AO22HSV2 U29 ( .A1(mux_bq[7]), .A2(n11), .B1(b_out[7]), .B2(n18), .Z(
        mux_b[7]) );
  LVT_AO22HSV4 U30 ( .A1(ti_7[0]), .A2(ctro), .B1(t_i_2_out[0]), .B2(n20), .Z(
        to_7[0]) );
  LVT_AO22HSV4 U31 ( .A1(ti_7[2]), .A2(ctro), .B1(t_i_2_out[2]), .B2(n20), .Z(
        to_7[2]) );
  LVT_AO22HSV4 U32 ( .A1(ti_7[4]), .A2(ctro), .B1(t_i_2_out[4]), .B2(n20), .Z(
        to_7[4]) );
  LVT_AO22HSV4 U33 ( .A1(ti_7[6]), .A2(ctro), .B1(t_i_2_out[6]), .B2(n20), .Z(
        to_7[6]) );
  LVT_INHSV2 U34 ( .I(rstn), .ZN(n15) );
endmodule


module regist_8bit_11 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_10 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_9 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_7 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_6 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_7 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV4 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV4 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV4 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_6 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_1bit_5 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_8 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_4 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_5 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module cell_3_99 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_13 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U3 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_XOR2HSV0 U5 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_12 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n2), .A3(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_11 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_10 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U3 ( .A1(n6), .A2(n5), .Z(n7) );
endmodule


module cell_4_9 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n2, n4;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_XNOR3HSV1 U2 ( .A1(n1), .A2(n4), .A3(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U3 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n1) );
endmodule


module cell_4_8 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n2), .A3(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_7 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n13) );
  LVT_NAND2HSV2 U2 ( .A1(n5), .A2(n6), .ZN(n14) );
  LVT_NAND2HSV2 U3 ( .A1(n1), .A2(n3), .ZN(n6) );
  LVT_INHSV2 U4 ( .I(n7), .ZN(n3) );
  LVT_INHSV2 U5 ( .I(n14), .ZN(n8) );
  LVT_NAND2HSV4 U6 ( .A1(n11), .A2(n10), .ZN(t_i_out) );
  LVT_CLKAND2HSV2 U7 ( .A1(b_in), .A2(a_in), .Z(n7) );
  LVT_XNOR2HSV1 U8 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n12) );
  LVT_CLKNHSV2 U9 ( .I(n13), .ZN(n1) );
  LVT_CLKNAND2HSV0 U10 ( .A1(n7), .A2(n13), .ZN(n5) );
  LVT_NAND2HSV2 U11 ( .A1(n14), .A2(n12), .ZN(n10) );
  LVT_NAND2HSV4 U12 ( .A1(n8), .A2(n9), .ZN(n11) );
  LVT_CLKNHSV2 U13 ( .I(n12), .ZN(n9) );
endmodule


module row_1_1 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_3_99 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_13 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(
        t_i_1_out[1]) );
  cell_4_12 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_11 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(
        t_i_1_out[3]) );
  cell_4_10 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(
        t_i_1_out[4]) );
  cell_4_9 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(t_i_1_out[5])
         );
  cell_4_8 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_7 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_13 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_98 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_97 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_96 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_95 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_94 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_93 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_XNOR2HSV1 U1 ( .A1(n6), .A2(n4), .ZN(t_i_out) );
  LVT_OAI21HSV2 U2 ( .A1(t_i_1_in), .A2(n5), .B(n2), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_NAND2HSV2 U5 ( .A1(n5), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_92 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;

  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n13) );
  LVT_CLKNAND2HSV2 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U3 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U4 ( .I(n13), .ZN(n2) );
  LVT_INHSV2SR U5 ( .I(n11), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(n11), .A2(n13), .ZN(n5) );
  LVT_CLKNAND2HSV1 U7 ( .A1(n7), .A2(n8), .ZN(n10) );
  LVT_CLKNHSV0P5 U8 ( .I(t_i_1_in), .ZN(n8) );
  LVT_NAND2HSV2 U9 ( .A1(n9), .A2(n10), .ZN(n11) );
  LVT_CLKNAND2HSV0 U10 ( .A1(n12), .A2(t_i_1_in), .ZN(n9) );
  LVT_INHSV2 U11 ( .I(n12), .ZN(n7) );
  LVT_NAND2HSV0 U12 ( .A1(b_in), .A2(a_in), .ZN(n12) );
endmodule


module row_other_13 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_13 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_98 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_97 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_96 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_95 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_94 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_93 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_92 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_12 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_91 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_90 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_89 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_88 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_87 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_86 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_85 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module row_other_12 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_12 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_91 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_90 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_89 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_88 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_87 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_86 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_85 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_11 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_84 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_83 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_82 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_81 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_80 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_79 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_78 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U4 ( .I(t_i_1_in), .ZN(n4) );
  LVT_NAND2HSV2 U5 ( .A1(n8), .A2(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV2 U6 ( .A1(n5), .A2(n6), .ZN(n7) );
  LVT_INHSV2 U7 ( .I(n8), .ZN(n2) );
  LVT_XNOR2HSV4 U8 ( .A1(n9), .A2(n7), .ZN(t_i_out) );
endmodule


module row_other_11 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_11 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_84 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_83 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_82 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_81 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_80 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_79 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_78 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_10 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_77 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_76 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_75 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_74 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_73 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_72 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_71 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV4 U1 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2SR U2 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV4 U5 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U6 ( .A1(n7), .A2(n9), .ZN(n5) );
  LVT_INHSV2 U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_10 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_10 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_77 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_76 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_75 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_74 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_73 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_72 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_71 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_9 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_70 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n10) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n11) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n12) );
  LVT_INHSV0P5 U4 ( .I(n12), .ZN(n6) );
  LVT_NAND2HSV0 U5 ( .A1(n7), .A2(n12), .ZN(n8) );
  LVT_CLKNAND2HSV0 U6 ( .A1(n6), .A2(n11), .ZN(n9) );
  LVT_NAND2HSV2 U7 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U8 ( .I(n10), .ZN(n4) );
  LVT_NAND2HSV2 U9 ( .A1(n8), .A2(n9), .ZN(t_i_out) );
  LVT_CLKNHSV1 U10 ( .I(n11), .ZN(n7) );
endmodule


module cell_3_69 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_68 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_67 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_66 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_65 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_64 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  LVT_NAND2HSV4 U1 ( .A1(n10), .A2(n11), .ZN(n13) );
  LVT_INHSV2SR U2 ( .I(n13), .ZN(n5) );
  LVT_CLKNAND2HSV1 U3 ( .A1(n12), .A2(n9), .ZN(n10) );
  LVT_CLKNHSV2 U4 ( .I(t_i_1_in), .ZN(n9) );
  LVT_CLKNAND2HSV3 U5 ( .A1(n4), .A2(n13), .ZN(n7) );
  LVT_CLKNAND2HSV3 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n14) );
  LVT_CLKNAND2HSV1 U7 ( .A1(n5), .A2(n14), .ZN(n6) );
  LVT_INHSV2 U8 ( .I(n14), .ZN(n4) );
  LVT_NAND2HSV1 U9 ( .A1(n8), .A2(t_i_1_in), .ZN(n11) );
  LVT_CLKNAND2HSV3 U10 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV2 U11 ( .I(n12), .ZN(n8) );
  LVT_NAND2HSV0 U12 ( .A1(b_in), .A2(a_in), .ZN(n12) );
endmodule


module row_other_9 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_9 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_70 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_69 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_68 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_67 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_66 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_65 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_64 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_8 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_63 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV2 U1 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_INHSV0P5SR U2 ( .I(n10), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(g_in), .A2(t_m_1_in), .ZN(n10) );
  LVT_NAND2HSV0P5 U5 ( .A1(n5), .A2(n10), .ZN(n6) );
  LVT_NAND2HSV0P5 U6 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_NAND2HSV2 U7 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV0SR U8 ( .I(n9), .ZN(n5) );
endmodule


module cell_3_62 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_61 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_60 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_59 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_58 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_AND2HSV0RD U1 ( .A1(b_in), .A2(a_in), .Z(n3) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV2 U3 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n3), .ZN(n4) );
endmodule


module cell_3_57 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV2 U1 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV0P5 U2 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV4 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNHSV4 U5 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_8 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_8 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_63 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_62 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_61 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_60 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_59 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_58 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_57 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_7 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_56 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INAND2HSV2 U2 ( .A1(n9), .B1(n8), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n7), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U5 ( .A1(n9), .A2(n4), .ZN(n5) );
  LVT_CLKNAND2HSV0 U6 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNHSV1 U7 ( .I(n8), .ZN(n4) );
endmodule


module cell_3_55 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_54 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_53 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_CLKNAND2HSV1 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U5 ( .I(n6), .ZN(n4) );
  LVT_XOR2HSV0 U6 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_3_52 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_51 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_50 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module row_other_7 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_7 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_56 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_55 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_54 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_53 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_52 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_51 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_50 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_1 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_1 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), .t_i_1_out(t0), 
        .t_i_2_out(t_i_2_out[6]) );
  row_other_13 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_12 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_11 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_10 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_9 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_8 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_7 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_7 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_6 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_7bit_4 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module PE_1 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   n24, l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17, n18, n19, n20, n21,
         n22, n23;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  LVT_AO22HSV0 U11 ( .A1(mux_bq[7]), .A2(n16), .B1(b_out[7]), .B2(n11), .Z(
        mux_b[7]) );
  LVT_AO22HSV0 U13 ( .A1(mux_bq[5]), .A2(n16), .B1(b_out[5]), .B2(n11), .Z(
        mux_b[5]) );
  LVT_AO22HSV0 U14 ( .A1(mux_bq[4]), .A2(n16), .B1(b_out[4]), .B2(n11), .Z(
        mux_b[4]) );
  LVT_AO22HSV0 U18 ( .A1(mux_bq[0]), .A2(n16), .B1(b_out[0]), .B2(n11), .Z(
        mux_b[0]) );
  regist_8bit_11 u0 ( .clk(clk), .rstn(n17), .in(a_in), .out(l_a) );
  regist_8bit_10 u1 ( .clk(clk), .rstn(n17), .in(b_in), .out(b_out) );
  regist_8bit_9 u2 ( .clk(clk), .rstn(n17), .in(g_in), .out(l_g) );
  regist_1bit_7 u3 ( .clk(clk), .rstn(n17), .in(ctr), .out(l_ctr) );
  regist_1bit_6 u4 ( .clk(clk), .rstn(n17), .in(n16), .out(ctro) );
  regist_7bit_7 u5 ( .clk(clk), .rstn(n17), .in(t_i_1_in), .out(l_t_i_1_in) );
  regist_7bit_6 u6 ( .clk(clk), .rstn(n17), .in(t_i_2_in), .out(l_t_i_2_in) );
  regist_1bit_5 u7 ( .clk(clk), .rstn(n17), .in(t_i_1_in_0), .out(l_t_i_1_in_0) );
  regist_8bit_8 u9 ( .clk(clk), .rstn(n17), .in(mux_b), .out(mux_bq) );
  regist_1bit_4 u10 ( .clk(clk), .rstn(n17), .in(n13), .out(ti_1) );
  regist_7bit_5 u11 ( .clk(clk), .rstn(n17), .in(to_7), .out(ti_7) );
  PE_core_1 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out({t_i_2_out[6], n24, t_i_2_out[4:0]}), 
        .t_i_1_out_0(t_i_1_out_0) );
  regist_8bit_7 u12 ( .clk(clk), .rstn(n17), .in(ao), .out(a_out) );
  regist_8bit_6 u13 ( .clk(clk), .rstn(n17), .in(go), .out(g_out) );
  regist_7bit_4 u14 ( .clk(clk), .rstn(n17), .in(to), .out(t_i_1_out) );
  LVT_CLKNAND2HSV8 U2 ( .A1(n8), .A2(n9), .ZN(to_7[2]) );
  LVT_INHSV0P5 U3 ( .I(l_ctr), .ZN(n21) );
  LVT_NOR2HSV2 U4 ( .A1(n22), .A2(n10), .ZN(c_t_i_1_in_0) );
  LVT_AO22HSV1 U5 ( .A1(mux_bq[2]), .A2(n16), .B1(b_out[2]), .B2(n10), .Z(
        mux_b[2]) );
  LVT_INHSV0SR U6 ( .I(n10), .ZN(n16) );
  LVT_AO22HSV1 U7 ( .A1(mux_bq[3]), .A2(n16), .B1(b_out[3]), .B2(n10), .Z(
        mux_b[3]) );
  LVT_AO22HSV1 U8 ( .A1(mux_bq[1]), .A2(n16), .B1(b_out[1]), .B2(n10), .Z(
        mux_b[1]) );
  LVT_AO22HSV1 U9 ( .A1(mux_bq[6]), .A2(n16), .B1(b_out[6]), .B2(n10), .Z(
        mux_b[6]) );
  LVT_CLKBUFHSV4 U10 ( .I(n21), .Z(n10) );
  LVT_INHSV2 U12 ( .I(ctro), .ZN(n23) );
  LVT_BUFHSV2 U15 ( .I(n21), .Z(n11) );
  LVT_NAND2HSV4 U16 ( .A1(ti_7[6]), .A2(ctro), .ZN(n6) );
  LVT_CLKNAND2HSV4 U17 ( .A1(t_i_2_out[6]), .A2(n23), .ZN(n7) );
  LVT_NAND2HSV8 U19 ( .A1(n6), .A2(n7), .ZN(to_7[6]) );
  LVT_NAND2HSV8 U20 ( .A1(ti_7[2]), .A2(ctro), .ZN(n8) );
  LVT_CLKNAND2HSV8 U21 ( .A1(t_i_2_out[2]), .A2(n23), .ZN(n9) );
  LVT_INHSV6 U22 ( .I(n18), .ZN(n17) );
  LVT_INHSV0SR U23 ( .I(to_1), .ZN(n12) );
  LVT_INHSV2 U24 ( .I(n12), .ZN(n13) );
  LVT_AOI21HSV2 U25 ( .A1(n20), .A2(n19), .B(n11), .ZN(\c_t_i_1_in[0] ) );
  LVT_NOR3HSV2 U26 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), .ZN(n20) );
  LVT_INHSV4SR U27 ( .I(l_t_i_1_in_0), .ZN(n22) );
  LVT_NOR4HSV12 U28 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(
        l_t_i_1_in[4]), .A4(l_t_i_1_in[3]), .ZN(n19) );
  LVT_INHSV0SR U29 ( .I(n24), .ZN(n14) );
  LVT_INHSV2 U30 ( .I(n14), .ZN(t_i_2_out[5]) );
  LVT_AO22HSV4 U31 ( .A1(ti_7[3]), .A2(ctro), .B1(t_i_2_out[3]), .B2(n23), .Z(
        to_7[3]) );
  LVT_AO22HSV4 U32 ( .A1(ti_7[5]), .A2(ctro), .B1(n24), .B2(n23), .Z(to_7[5])
         );
  LVT_AO22HSV4 U33 ( .A1(ti_7[0]), .A2(ctro), .B1(t_i_2_out[0]), .B2(n23), .Z(
        to_7[0]) );
  LVT_AO22HSV4 U34 ( .A1(ti_7[1]), .A2(ctro), .B1(t_i_2_out[1]), .B2(n23), .Z(
        to_7[1]) );
  LVT_AO22HSV4 U35 ( .A1(ti_7[4]), .A2(ctro), .B1(t_i_2_out[4]), .B2(n23), .Z(
        to_7[4]) );
  LVT_MOAI22HSV4 U36 ( .A1(l_ctr), .A2(n22), .B1(l_ctr), .B2(ti_1), .ZN(to_1)
         );
  LVT_INHSV2 U37 ( .I(rstn), .ZN(n18) );
endmodule


module regist_8bit_5 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_4 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_8bit_3 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_3 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_2 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_3 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV4 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV4 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV4 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV4 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_7bit_2 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
endmodule


module regist_1bit_1 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_8bit_2 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n2) );
endmodule


module regist_1bit_0 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_7bit_1 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module cell_3_49 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_6 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_5 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_4 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_3 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_XOR3HSV1 U2 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
endmodule


module cell_4_2 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV2 U1 ( .A1(n5), .A2(n2), .A3(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_1 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n2, n4;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR3HSV2 U1 ( .A1(n1), .A2(n2), .A3(n4), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_XNOR2HSV1 U3 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n1) );
endmodule


module cell_4_0 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10, n11;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n10) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV1 U2 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_CLKXOR2HSV2 U3 ( .A1(n9), .A2(n10), .Z(n11) );
  LVT_XNOR2HSV1 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n8) );
  LVT_INHSV2SR U6 ( .I(n11), .ZN(n5) );
  LVT_NAND2HSV2 U7 ( .A1(n1), .A2(n5), .ZN(n7) );
  LVT_INHSV2 U8 ( .I(n8), .ZN(n1) );
  LVT_CLKNAND2HSV0 U9 ( .A1(n8), .A2(n11), .ZN(n6) );
endmodule


module row_1_0 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_3_49 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_6 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(
        t_i_1_out[1]) );
  cell_4_5 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(
        t_i_1_out[2]) );
  cell_4_4 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(
        t_i_1_out[3]) );
  cell_4_3 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(
        t_i_1_out[4]) );
  cell_4_2 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(
        t_i_1_out[5]) );
  cell_4_1 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(
        t_i_1_out[6]) );
  cell_4_0 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_6 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_48 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_47 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_46 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n8), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(n8), .A2(n4), .ZN(n5) );
  LVT_CLKNHSV0 U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_45 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_44 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_43 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_42 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV0 U2 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2 U4 ( .I(n9), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV4 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U7 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNAND2HSV3 U8 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
endmodule


module row_other_6 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_6 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_48 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_47 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_46 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_45 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_44 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_43 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_42 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_5 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_41 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4;

  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n4) );
  LVT_CLKAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .Z(n2) );
  LVT_XOR2HSV4 U3 ( .A1(n2), .A2(t_i_1_in), .Z(n3) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(n3), .ZN(t_i_out) );
endmodule


module cell_3_40 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_39 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_38 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_37 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(g_in), .A2(t_m_1_in), .ZN(n6) );
endmodule


module cell_3_36 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_35 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV2 U2 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV3SR U5 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV4 U6 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_INHSV2 U7 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV1 U8 ( .A1(n9), .A2(n7), .ZN(n5) );
endmodule


module row_other_5 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_5 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_41 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_40 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_39 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_38 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_37 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_36 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_35 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_4 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(n3), .Z(t_i_out) );
endmodule


module cell_3_34 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_33 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_32 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_31 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_30 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_29 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_NAND2HSV2 U1 ( .A1(n6), .A2(t_i_1_in), .ZN(n7) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(n9), .B(n5), .ZN(t_i_out) );
  LVT_OAI21HSV2 U3 ( .A1(n6), .A2(t_i_1_in), .B(n7), .ZN(n9) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(n9), .ZN(n5) );
  LVT_INHSV2 U6 ( .I(n10), .ZN(n4) );
  LVT_CLKNHSV0P5 U7 ( .I(n8), .ZN(n6) );
  LVT_NAND2HSV0 U8 ( .A1(b_in), .A2(a_in), .ZN(n8) );
endmodule


module cell_3_28 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV2 U1 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_NAND2HSV2 U5 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV4 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV3 U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_4 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_4 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_34 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_33 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_32 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_31 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_30 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_29 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_28 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_3 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_XOR2HSV0 U2 ( .A1(n3), .A2(n4), .Z(t_i_out) );
endmodule


module cell_3_27 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_26 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_25 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_24 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_23 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_22 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_21 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XNOR2HSV1 U1 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
  LVT_INHSV2 U2 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV3 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV0 U5 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV3SR U6 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV4 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U8 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
endmodule


module row_other_3 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_3 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_27 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_26 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_25 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_24 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_23 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_22 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_21 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_2 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_20 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_19 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_18 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_17 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_16 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_15 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_14 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2SR U4 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV0P5 U5 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV4 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV2SR U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_2 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_2 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_20 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_19 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_18 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_17 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_16 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_15 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_14 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_1 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_13 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_12 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_11 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_10 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_9 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_8 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_7 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV2 U2 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV1 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV4 U5 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV4 U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_1 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_1 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_13 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_12 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_11 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_10 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_9 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_8 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_7 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_0 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4, n5, n6;

  LVT_OAI21HSV2 U1 ( .A1(n3), .A2(n5), .B(n4), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U3 ( .A1(n3), .A2(n5), .ZN(n4) );
  LVT_INHSV0SR U4 ( .I(n6), .ZN(n3) );
  LVT_NAND2HSV0P5 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_6 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_5 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_INHSV2SR U5 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0P5 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_4 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_3 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_INHSV1SR U5 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0P5 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_2 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_1 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_0 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U2 ( .A1(g_in), .A2(t_m_1_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module row_other_0 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [7:0] a_in;
  input [7:0] g_in;
  input [6:0] t_i_1_in;
  output [6:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_0 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_6 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_0 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_0 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [7:0] t_m_1_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;

  wire   [6:0] t0;
  wire   [6:0] t1;
  wire   [6:0] t2;
  wire   [6:0] t3;
  wire   [6:0] t4;
  wire   [6:0] t5;
  wire   [6:0] t6;
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_0 u0 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[7]), .t_m_1_in(t_m_1_in[7]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), .t_i_1_out(t0), 
        .t_i_2_out(t_i_2_out[6]) );
  row_other_6 u1 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[6]), .t_m_1_in(
        t_m_1_in[6]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[5])
         );
  row_other_5 u2 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[5]), .t_m_1_in(
        t_m_1_in[5]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[4])
         );
  row_other_4 u3 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[4]), .t_m_1_in(
        t_m_1_in[4]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[3])
         );
  row_other_3 u4 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[3]), .t_m_1_in(
        t_m_1_in[3]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[2])
         );
  row_other_2 u5 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[2]), .t_m_1_in(
        t_m_1_in[2]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[1])
         );
  row_other_1 u6 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[1]), .t_m_1_in(
        t_m_1_in[1]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[0])
         );
  row_other_0 u7 ( .a_in(a_in), .g_in(g_in), .b_in(b_in[0]), .t_m_1_in(
        t_m_1_in[0]), .t_i_1_in(t6), .t_i_1_out(t_i_1_out), .t_i_2_out(
        t_i_1_out_0) );
endmodule


module regist_8bit_1 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_8bit_0 ( clk, rstn, in, out );
  input [7:0] in;
  output [7:0] out;
  input clk, rstn;


  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module regist_7bit_0 ( clk, rstn, in, out );
  input [6:0] in;
  output [6:0] out;
  input clk, rstn;


  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
endmodule


module PE_0 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  input [6:0] t_i_1_in;
  input [6:0] t_i_2_in;
  output [7:0] a_out;
  output [7:0] g_out;
  output [7:0] b_out;
  output [6:0] t_i_1_out;
  output [6:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23;
  wire   [7:0] l_a;
  wire   [7:0] l_g;
  wire   [6:0] l_t_i_1_in;
  wire   [6:0] l_t_i_2_in;
  wire   [7:0] mux_b;
  wire   [7:0] mux_bq;
  wire   [6:0] to_7;
  wire   [6:0] ti_7;
  wire   [7:0] ao;
  wire   [7:0] go;
  wire   [6:0] to;

  LVT_NOR3HSV0 U24 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[2]), .A3(l_t_i_1_in[1]), .ZN(n20) );
  regist_8bit_5 u0 ( .clk(clk), .rstn(n17), .in(a_in), .out(l_a) );
  regist_8bit_4 u1 ( .clk(clk), .rstn(n17), .in(b_in), .out(b_out) );
  regist_8bit_3 u2 ( .clk(clk), .rstn(n17), .in(g_in), .out(l_g) );
  regist_1bit_3 u3 ( .clk(clk), .rstn(n17), .in(ctr), .out(l_ctr) );
  regist_1bit_2 u4 ( .clk(clk), .rstn(n17), .in(n16), .out(ctro) );
  regist_7bit_3 u5 ( .clk(clk), .rstn(n17), .in(t_i_1_in), .out(l_t_i_1_in) );
  regist_7bit_2 u6 ( .clk(clk), .rstn(n17), .in(t_i_2_in), .out(l_t_i_2_in) );
  regist_1bit_1 u7 ( .clk(clk), .rstn(n17), .in(t_i_1_in_0), .out(l_t_i_1_in_0) );
  regist_8bit_2 u9 ( .clk(clk), .rstn(n17), .in(mux_b), .out(mux_bq) );
  regist_1bit_0 u10 ( .clk(clk), .rstn(n17), .in(n15), .out(ti_1) );
  regist_7bit_1 u11 ( .clk(clk), .rstn(n17), .in(to_7), .out(ti_7) );
  PE_core_0 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out(t_i_2_out), .t_i_1_out_0(t_i_1_out_0)
         );
  regist_8bit_1 u12 ( .clk(clk), .rstn(n17), .in(ao), .out(a_out) );
  regist_8bit_0 u13 ( .clk(clk), .rstn(n17), .in(go), .out(g_out) );
  regist_7bit_0 u14 ( .clk(clk), .rstn(n17), .in(to), .out(t_i_1_out) );
  LVT_NAND2HSV8 U2 ( .A1(n8), .A2(n9), .ZN(to_7[0]) );
  LVT_INHSV4SR U3 ( .I(n12), .ZN(n13) );
  LVT_CLKNAND2HSV4 U4 ( .A1(t_i_2_out[0]), .A2(n23), .ZN(n9) );
  LVT_CLKNAND2HSV4 U5 ( .A1(n6), .A2(n7), .ZN(to_7[6]) );
  LVT_INHSV2 U6 ( .I(n21), .ZN(n12) );
  LVT_INHSV2 U7 ( .I(ctro), .ZN(n23) );
  LVT_NOR2HSV1 U8 ( .A1(n22), .A2(n13), .ZN(c_t_i_1_in_0) );
  LVT_NAND2HSV2 U9 ( .A1(ti_7[6]), .A2(ctro), .ZN(n6) );
  LVT_CLKNAND2HSV3 U10 ( .A1(t_i_2_out[6]), .A2(n23), .ZN(n7) );
  LVT_CLKNAND2HSV1 U11 ( .A1(ti_7[0]), .A2(ctro), .ZN(n8) );
  LVT_CLKNAND2HSV8 U12 ( .A1(ti_7[4]), .A2(ctro), .ZN(n10) );
  LVT_CLKNAND2HSV8 U13 ( .A1(t_i_2_out[4]), .A2(n23), .ZN(n11) );
  LVT_NAND2HSV8 U14 ( .A1(n10), .A2(n11), .ZN(to_7[4]) );
  LVT_INHSV0SR U15 ( .I(l_ctr), .ZN(n21) );
  LVT_INHSV6 U16 ( .I(n18), .ZN(n17) );
  LVT_INHSV0SR U17 ( .I(to_1), .ZN(n14) );
  LVT_INHSV2 U18 ( .I(n14), .ZN(n15) );
  LVT_INHSV2 U19 ( .I(l_t_i_1_in_0), .ZN(n22) );
  LVT_BUFHSV2RT U20 ( .I(l_ctr), .Z(n16) );
  LVT_NOR4HSV12 U21 ( .A1(l_t_i_1_in[6]), .A2(l_t_i_1_in[5]), .A3(
        l_t_i_1_in[4]), .A4(l_t_i_1_in[3]), .ZN(n19) );
  LVT_AOI21HSV0 U22 ( .A1(n20), .A2(n19), .B(n13), .ZN(\c_t_i_1_in[0] ) );
  LVT_AO22HSV2 U23 ( .A1(mux_bq[1]), .A2(n16), .B1(b_out[1]), .B2(n13), .Z(
        mux_b[1]) );
  LVT_AO22HSV2 U25 ( .A1(mux_bq[2]), .A2(n16), .B1(b_out[2]), .B2(n13), .Z(
        mux_b[2]) );
  LVT_AO22HSV2 U26 ( .A1(mux_bq[3]), .A2(n16), .B1(b_out[3]), .B2(n13), .Z(
        mux_b[3]) );
  LVT_AO22HSV2 U27 ( .A1(mux_bq[4]), .A2(n16), .B1(b_out[4]), .B2(n13), .Z(
        mux_b[4]) );
  LVT_AO22HSV2 U28 ( .A1(mux_bq[0]), .A2(n16), .B1(b_out[0]), .B2(n13), .Z(
        mux_b[0]) );
  LVT_AO22HSV2 U29 ( .A1(mux_bq[7]), .A2(l_ctr), .B1(b_out[7]), .B2(n13), .Z(
        mux_b[7]) );
  LVT_AO22HSV4 U30 ( .A1(ti_7[5]), .A2(ctro), .B1(t_i_2_out[5]), .B2(n23), .Z(
        to_7[5]) );
  LVT_AO22HSV2 U31 ( .A1(mux_bq[6]), .A2(n16), .B1(b_out[6]), .B2(n13), .Z(
        mux_b[6]) );
  LVT_AO22HSV2 U32 ( .A1(mux_bq[5]), .A2(n16), .B1(b_out[5]), .B2(n13), .Z(
        mux_b[5]) );
  LVT_AO22HSV4 U33 ( .A1(ti_7[1]), .A2(ctro), .B1(t_i_2_out[1]), .B2(n23), .Z(
        to_7[1]) );
  LVT_AO22HSV4 U34 ( .A1(ti_7[2]), .A2(ctro), .B1(t_i_2_out[2]), .B2(n23), .Z(
        to_7[2]) );
  LVT_AO22HSV4 U35 ( .A1(ti_7[3]), .A2(ctro), .B1(t_i_2_out[3]), .B2(n23), .Z(
        to_7[3]) );
  LVT_INHSV2 U36 ( .I(rstn), .ZN(n18) );
  LVT_MOAI22HSV4 U37 ( .A1(l_ctr), .A2(n22), .B1(ti_1), .B2(l_ctr), .ZN(to_1)
         );
endmodule


module regist_1bit_84 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module top ( clk, rstn, ctr, a_in, g_in, b_in, po, ctro );
  input [7:0] a_in;
  input [7:0] g_in;
  input [7:0] b_in;
  output [7:0] po;
  input clk, rstn, ctr;
  output ctro;
  wire   po1, ctro1, po2, ctro2, po3, ctro3, po4, ctro4, po5, ctro5, po6,
         ctro6, po7, ctro7, po8, ctro8, po9, ctro9, po10, ctro10, po11, ctro11,
         po12, ctro12, po13, ctro13, po14, ctro14, po15, ctro15, po16, ctro16,
         po17, ctro17, po18, ctro18, po19, ctro19, po20, ctro20, po21, n1, n2,
         n3, n4, n5, n6, n7;
  wire   [7:0] ao1;
  wire   [7:0] go1;
  wire   [7:0] bo1;
  wire   [6:0] poh1;
  wire   [6:0] pov1;
  wire   [7:0] ao2;
  wire   [7:0] go2;
  wire   [7:0] bo2;
  wire   [6:0] poh2;
  wire   [6:0] pov2;
  wire   [7:0] ao3;
  wire   [7:0] go3;
  wire   [7:0] bo3;
  wire   [6:0] poh3;
  wire   [6:0] pov3;
  wire   [7:0] ao4;
  wire   [7:0] go4;
  wire   [7:0] bo4;
  wire   [6:0] poh4;
  wire   [6:0] pov4;
  wire   [7:0] ao5;
  wire   [7:0] go5;
  wire   [7:0] bo5;
  wire   [6:0] poh5;
  wire   [6:0] pov5;
  wire   [7:0] ao6;
  wire   [7:0] go6;
  wire   [7:0] bo6;
  wire   [6:0] poh6;
  wire   [6:0] pov6;
  wire   [7:0] ao7;
  wire   [7:0] go7;
  wire   [7:0] bo7;
  wire   [6:0] poh7;
  wire   [6:0] pov7;
  wire   [7:0] ao8;
  wire   [7:0] go8;
  wire   [7:0] bo8;
  wire   [6:0] poh8;
  wire   [6:0] pov8;
  wire   [7:0] ao9;
  wire   [7:0] go9;
  wire   [7:0] bo9;
  wire   [6:0] poh9;
  wire   [6:0] pov9;
  wire   [7:0] ao10;
  wire   [7:0] go10;
  wire   [7:0] bo10;
  wire   [6:0] poh10;
  wire   [6:0] pov10;
  wire   [7:0] ao11;
  wire   [7:0] go11;
  wire   [7:0] bo11;
  wire   [6:0] poh11;
  wire   [6:0] pov11;
  wire   [7:0] ao12;
  wire   [7:0] go12;
  wire   [7:0] bo12;
  wire   [6:0] poh12;
  wire   [6:0] pov12;
  wire   [7:0] ao13;
  wire   [7:0] go13;
  wire   [7:0] bo13;
  wire   [6:0] poh13;
  wire   [6:0] pov13;
  wire   [7:0] ao14;
  wire   [7:0] go14;
  wire   [7:0] bo14;
  wire   [6:0] poh14;
  wire   [6:0] pov14;
  wire   [7:0] ao15;
  wire   [7:0] go15;
  wire   [7:0] bo15;
  wire   [6:0] poh15;
  wire   [6:0] pov15;
  wire   [7:0] ao16;
  wire   [7:0] go16;
  wire   [7:0] bo16;
  wire   [6:0] poh16;
  wire   [6:0] pov16;
  wire   [7:0] ao17;
  wire   [7:0] go17;
  wire   [7:0] bo17;
  wire   [6:0] poh17;
  wire   [6:0] pov17;
  wire   [7:0] ao18;
  wire   [7:0] go18;
  wire   [7:0] bo18;
  wire   [6:0] poh18;
  wire   [6:0] pov18;
  wire   [7:0] ao19;
  wire   [7:0] go19;
  wire   [7:0] bo19;
  wire   [6:0] poh19;
  wire   [6:0] pov19;
  wire   [7:0] ao20;
  wire   [7:0] go20;
  wire   [7:0] bo20;
  wire   [6:0] poh20;
  wire   [6:0] pov20;
  wire   [6:0] poh21;
  wire   [6:0] pov21;

  PE_20 pe0 ( .clk(clk), .rstn(rstn), .ctr(ctr), .a_in(a_in), .g_in(g_in), 
        .b_in(b_in), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .t_i_1_in_0(1'b0), .t_i_2_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a_out(ao1), .g_out(go1), .b_out(bo1), .t_i_1_out(poh1), .t_i_2_out(pov1), 
        .t_i_1_out_0(po1), .ctro(ctro1) );
  PE_19 pe1 ( .clk(clk), .rstn(rstn), .ctr(ctro1), .a_in(ao1), .g_in(go1), 
        .b_in(bo1), .t_i_1_in(poh1), .t_i_1_in_0(po1), .t_i_2_in(pov1), 
        .a_out(ao2), .g_out(go2), .b_out(bo2), .t_i_1_out(poh2), .t_i_2_out(
        pov2), .t_i_1_out_0(po2), .ctro(ctro2) );
  PE_18 pe2 ( .clk(clk), .rstn(rstn), .ctr(ctro2), .a_in(ao2), .g_in(go2), 
        .b_in(bo2), .t_i_1_in(poh2), .t_i_1_in_0(po2), .t_i_2_in(pov2), 
        .a_out(ao3), .g_out(go3), .b_out(bo3), .t_i_1_out(poh3), .t_i_2_out(
        pov3), .t_i_1_out_0(po3), .ctro(ctro3) );
  PE_17 pe3 ( .clk(clk), .rstn(rstn), .ctr(ctro3), .a_in(ao3), .g_in(go3), 
        .b_in(bo3), .t_i_1_in(poh3), .t_i_1_in_0(po3), .t_i_2_in(pov3), 
        .a_out(ao4), .g_out(go4), .b_out(bo4), .t_i_1_out(poh4), .t_i_2_out(
        pov4), .t_i_1_out_0(po4), .ctro(ctro4) );
  PE_16 pe4 ( .clk(clk), .rstn(rstn), .ctr(ctro4), .a_in(ao4), .g_in(go4), 
        .b_in(bo4), .t_i_1_in(poh4), .t_i_1_in_0(po4), .t_i_2_in(pov4), 
        .a_out(ao5), .g_out(go5), .b_out(bo5), .t_i_1_out(poh5), .t_i_2_out(
        pov5), .t_i_1_out_0(po5), .ctro(ctro5) );
  PE_15 pe5 ( .clk(clk), .rstn(rstn), .ctr(ctro5), .a_in(ao5), .g_in(go5), 
        .b_in(bo5), .t_i_1_in(poh5), .t_i_1_in_0(po5), .t_i_2_in(pov5), 
        .a_out(ao6), .g_out(go6), .b_out(bo6), .t_i_1_out(poh6), .t_i_2_out(
        pov6), .t_i_1_out_0(po6), .ctro(ctro6) );
  PE_14 pe6 ( .clk(clk), .rstn(rstn), .ctr(ctro6), .a_in(ao6), .g_in(go6), 
        .b_in(bo6), .t_i_1_in(poh6), .t_i_1_in_0(po6), .t_i_2_in(pov6), 
        .a_out(ao7), .g_out(go7), .b_out(bo7), .t_i_1_out(poh7), .t_i_2_out(
        pov7), .t_i_1_out_0(po7), .ctro(ctro7) );
  PE_13 pe7 ( .clk(clk), .rstn(rstn), .ctr(ctro7), .a_in(ao7), .g_in(go7), 
        .b_in(bo7), .t_i_1_in(poh7), .t_i_1_in_0(po7), .t_i_2_in(pov7), 
        .a_out(ao8), .g_out(go8), .b_out(bo8), .t_i_1_out(poh8), .t_i_2_out(
        pov8), .t_i_1_out_0(po8), .ctro(ctro8) );
  PE_12 pe8 ( .clk(clk), .rstn(rstn), .ctr(ctro8), .a_in(ao8), .g_in(go8), 
        .b_in(bo8), .t_i_1_in(poh8), .t_i_1_in_0(po8), .t_i_2_in(pov8), 
        .a_out(ao9), .g_out(go9), .b_out(bo9), .t_i_1_out(poh9), .t_i_2_out(
        pov9), .t_i_1_out_0(po9), .ctro(ctro9) );
  PE_11 pe9 ( .clk(clk), .rstn(rstn), .ctr(ctro9), .a_in(ao9), .g_in(go9), 
        .b_in(bo9), .t_i_1_in(poh9), .t_i_1_in_0(po9), .t_i_2_in(pov9), 
        .a_out(ao10), .g_out(go10), .b_out(bo10), .t_i_1_out(poh10), 
        .t_i_2_out(pov10), .t_i_1_out_0(po10), .ctro(ctro10) );
  PE_10 pe10 ( .clk(clk), .rstn(rstn), .ctr(ctro10), .a_in(ao10), .g_in(go10), 
        .b_in(bo10), .t_i_1_in(poh10), .t_i_1_in_0(po10), .t_i_2_in(pov10), 
        .a_out(ao11), .g_out(go11), .b_out(bo11), .t_i_1_out(poh11), 
        .t_i_2_out(pov11), .t_i_1_out_0(po11), .ctro(ctro11) );
  PE_9 pe11 ( .clk(clk), .rstn(rstn), .ctr(ctro11), .a_in(ao11), .g_in(go11), 
        .b_in(bo11), .t_i_1_in(poh11), .t_i_1_in_0(po11), .t_i_2_in(pov11), 
        .a_out(ao12), .g_out(go12), .b_out(bo12), .t_i_1_out(poh12), 
        .t_i_2_out(pov12), .t_i_1_out_0(po12), .ctro(ctro12) );
  PE_8 pe12 ( .clk(clk), .rstn(rstn), .ctr(ctro12), .a_in(ao12), .g_in(go12), 
        .b_in(bo12), .t_i_1_in(poh12), .t_i_1_in_0(po12), .t_i_2_in(pov12), 
        .a_out(ao13), .g_out(go13), .b_out(bo13), .t_i_1_out(poh13), 
        .t_i_2_out(pov13), .t_i_1_out_0(po13), .ctro(ctro13) );
  PE_7 pe13 ( .clk(clk), .rstn(rstn), .ctr(ctro13), .a_in(ao13), .g_in(go13), 
        .b_in(bo13), .t_i_1_in(poh13), .t_i_1_in_0(po13), .t_i_2_in(pov13), 
        .a_out(ao14), .g_out(go14), .b_out(bo14), .t_i_1_out(poh14), 
        .t_i_2_out(pov14), .t_i_1_out_0(po14), .ctro(ctro14) );
  PE_6 pe14 ( .clk(clk), .rstn(rstn), .ctr(ctro14), .a_in(ao14), .g_in(go14), 
        .b_in(bo14), .t_i_1_in(poh14), .t_i_1_in_0(po14), .t_i_2_in(pov14), 
        .a_out(ao15), .g_out(go15), .b_out(bo15), .t_i_1_out(poh15), 
        .t_i_2_out(pov15), .t_i_1_out_0(po15), .ctro(ctro15) );
  PE_5 pe15 ( .clk(clk), .rstn(rstn), .ctr(ctro15), .a_in(ao15), .g_in(go15), 
        .b_in(bo15), .t_i_1_in(poh15), .t_i_1_in_0(po15), .t_i_2_in(pov15), 
        .a_out(ao16), .g_out(go16), .b_out(bo16), .t_i_1_out(poh16), 
        .t_i_2_out(pov16), .t_i_1_out_0(po16), .ctro(ctro16) );
  PE_4 pe16 ( .clk(clk), .rstn(rstn), .ctr(ctro16), .a_in(ao16), .g_in(go16), 
        .b_in(bo16), .t_i_1_in(poh16), .t_i_1_in_0(po16), .t_i_2_in(pov16), 
        .a_out(ao17), .g_out(go17), .b_out(bo17), .t_i_1_out(poh17), 
        .t_i_2_out(pov17), .t_i_1_out_0(po17), .ctro(ctro17) );
  PE_3 pe17 ( .clk(clk), .rstn(rstn), .ctr(ctro17), .a_in(ao17), .g_in(go17), 
        .b_in(bo17), .t_i_1_in(poh17), .t_i_1_in_0(po17), .t_i_2_in(pov17), 
        .a_out(ao18), .g_out(go18), .b_out(bo18), .t_i_1_out(poh18), 
        .t_i_2_out(pov18), .t_i_1_out_0(po18), .ctro(ctro18) );
  PE_2 pe18 ( .clk(clk), .rstn(rstn), .ctr(ctro18), .a_in(ao18), .g_in(go18), 
        .b_in(bo18), .t_i_1_in(poh18), .t_i_1_in_0(po18), .t_i_2_in(pov18), 
        .a_out(ao19), .g_out(go19), .b_out(bo19), .t_i_1_out(poh19), 
        .t_i_2_out(pov19), .t_i_1_out_0(po19), .ctro(ctro19) );
  PE_1 pe19 ( .clk(clk), .rstn(rstn), .ctr(ctro19), .a_in(ao19), .g_in(go19), 
        .b_in(bo19), .t_i_1_in(poh19), .t_i_1_in_0(po19), .t_i_2_in(pov19), 
        .a_out(ao20), .g_out(go20), .b_out(bo20), .t_i_1_out(poh20), 
        .t_i_2_out(pov20), .t_i_1_out_0(po20), .ctro(ctro20) );
  PE_0 pe20 ( .clk(clk), .rstn(rstn), .ctr(ctro20), .a_in(ao20), .g_in(go20), 
        .b_in(bo20), .t_i_1_in(poh20), .t_i_1_in_0(po20), .t_i_2_in(pov20), 
        .a_out(), .g_out(), .b_out(), .t_i_1_out(poh21), .t_i_2_out(pov21), 
        .t_i_1_out_0(po21), .ctro(ctro) );
  regist_1bit_84 pe21 ( .clk(clk), .rstn(rstn), .in(po21), .out(po[7]) );
  LVT_XOR2HSV0 U2 ( .A1(poh21[0]), .A2(n6), .Z(po[0]) );
  LVT_XOR2HSV0 U3 ( .A1(poh21[1]), .A2(n5), .Z(po[1]) );
  LVT_XOR2HSV0 U4 ( .A1(poh21[2]), .A2(n4), .Z(po[2]) );
  LVT_AND2HSV0RD U5 ( .A1(pov21[0]), .A2(ctro), .Z(n6) );
  LVT_AND2HSV0RD U6 ( .A1(pov21[1]), .A2(ctro), .Z(n5) );
  LVT_AND2HSV0RD U7 ( .A1(pov21[2]), .A2(ctro), .Z(n4) );
  LVT_XOR2HSV0 U8 ( .A1(poh21[3]), .A2(n3), .Z(po[3]) );
  LVT_AND2HSV0RD U9 ( .A1(pov21[3]), .A2(ctro), .Z(n3) );
  LVT_XOR2HSV0 U10 ( .A1(poh21[4]), .A2(n2), .Z(po[4]) );
  LVT_AND2HSV0RD U11 ( .A1(pov21[4]), .A2(ctro), .Z(n2) );
  LVT_XOR2HSV0 U12 ( .A1(poh21[5]), .A2(n1), .Z(po[5]) );
  LVT_AND2HSV0RD U13 ( .A1(pov21[5]), .A2(ctro), .Z(n1) );
  LVT_XNOR2HSV1 U14 ( .A1(poh21[6]), .A2(n7), .ZN(po[6]) );
  LVT_NAND2HSV0 U15 ( .A1(pov21[6]), .A2(ctro), .ZN(n7) );
endmodule

