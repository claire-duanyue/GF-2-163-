
module regist_32bit_35 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3, n4;

  LVT_DRNQHSV4 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV4 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV4 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV4 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV4 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV4 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV4 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n3), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n3), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n3), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n3), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n3), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n3), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n3), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n3), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_INHSV2 U3 ( .I(n4), .ZN(n2) );
  LVT_INHSV2 U4 ( .I(n4), .ZN(n1) );
  LVT_INHSV2 U5 ( .I(rstn), .ZN(n4) );
  LVT_INHSV2 U6 ( .I(n4), .ZN(n3) );
endmodule


module regist_32bit_34 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV2 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_32bit_33 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV4 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV4 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV4 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV4 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV4 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n2), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(rstn), .Q(out[19])
         );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(rstn), .Q(out[18])
         );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(rstn), .Q(out[17])
         );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(rstn), .Q(out[16])
         );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(rstn), .Q(out[15])
         );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(rstn), .Q(out[14])
         );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(rstn), .Q(out[13])
         );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n2), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n2), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n2), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_INHSV2 U3 ( .I(n3), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n2) );
endmodule


module regist_1bit_23 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_22 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_31bit_23 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n2), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n2), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n2), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n2), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n2), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n1), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n1), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n1), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n1), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n1), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n1), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n2), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n2), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n2), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n3), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n2) );
endmodule


module regist_31bit_22 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n2), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n2), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n2), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n2), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n2), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n2), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n1), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n1), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n1), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n1), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n1), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n1), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n2), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n2), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n3), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n2) );
endmodule


module regist_1bit_21 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_32bit_32 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n6, n1, n3, n4, n5;

  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n4), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n4), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n4), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n3), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n4), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n3), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n4), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n3), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n4), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n3), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n3), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n4), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n4), .Q(n6) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n4), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n4), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n4), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n3), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n3), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n3), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n3), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n3), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n3), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n3), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n3), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n3), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n3), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n3), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n4), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n4), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n4), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n4), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n4), .Q(out[12]) );
  LVT_INHSV8SR U3 ( .I(n1), .ZN(out[31]) );
  LVT_INHSV2 U4 ( .I(n6), .ZN(n1) );
  LVT_INHSV2 U5 ( .I(n5), .ZN(n3) );
  LVT_INHSV2 U6 ( .I(rstn), .ZN(n5) );
  LVT_INHSV2 U7 ( .I(n5), .ZN(n4) );
endmodule


module regist_1bit_20 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_31bit_21 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(rstn), .Q(out[30])
         );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n2), .Q(out[28]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(rstn), .Q(out[27])
         );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n2), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(rstn), .Q(out[24])
         );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n2), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n2), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n1) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n2) );
endmodule


module cell_3_5771 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n1, n2, n3;

  LVT_XOR2HSV0 U1 ( .A1(n1), .A2(n2), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n3), .A2(t_i_1_in), .Z(n2) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n1) );
endmodule


module cell_4_185 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n2, n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n1), .A2(n2), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n3), .A2(n4), .Z(n2) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n3) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n1) );
endmodule


module cell_4_184 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_183 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_182 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_181 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_180 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_179 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_178 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_177 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_176 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_175 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_174 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_173 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_172 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_171 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_170 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_169 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_168 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_167 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_NAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_4_166 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_4_165 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_4_164 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_163 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_4_162 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_161 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_160 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_159 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U3 ( .A1(n6), .A2(n5), .Z(n7) );
endmodule


module cell_4_158 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_157 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_XOR3HSV1 U2 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
endmodule


module cell_4_156 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n5, n6, n7, n8, n9, n10, n11;

  LVT_NAND2HSV2 U1 ( .A1(n2), .A2(n5), .ZN(n7) );
  LVT_INHSV1SR U2 ( .I(n10), .ZN(n2) );
  LVT_CLKNHSV2 U3 ( .I(n9), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n8), .A2(n11), .ZN(t_i_out) );
  LVT_NAND2HSV0 U5 ( .A1(n10), .A2(n9), .ZN(n6) );
  LVT_NAND2HSV1 U6 ( .A1(b_in), .A2(a_in), .ZN(n10) );
  LVT_NAND2HSV2 U7 ( .A1(n6), .A2(n7), .ZN(n8) );
  LVT_XOR2HSV0 U8 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n11) );
  LVT_CLKNAND2HSV2 U9 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
endmodule


module cell_4_155 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  LVT_NAND2HSV4 U1 ( .A1(n1), .A2(n5), .ZN(n6) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV2SR U3 ( .I(n15), .ZN(n1) );
  LVT_INHSV0P5SR U4 ( .I(n12), .ZN(n5) );
  LVT_XNOR2HSV4 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n12) );
  LVT_CLKNAND2HSV2 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n13) );
  LVT_INHSV2 U7 ( .I(n13), .ZN(n9) );
  LVT_NAND2HSV2 U8 ( .A1(n8), .A2(n13), .ZN(n11) );
  LVT_INHSV1SR U9 ( .I(n14), .ZN(n8) );
  LVT_NAND2HSV2 U10 ( .A1(b_in), .A2(a_in), .ZN(n14) );
  LVT_CLKNAND2HSV1 U11 ( .A1(n9), .A2(n14), .ZN(n10) );
  LVT_NAND2HSV2 U12 ( .A1(n10), .A2(n11), .ZN(n15) );
  LVT_NAND2HSV0P5 U13 ( .A1(n15), .A2(n12), .ZN(n7) );
endmodule


module row_1_5 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [31:0] t_i_1_in;
  input [30:0] t_i_2_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_3_5771 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_185 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(t_i_1_out[1])
         );
  cell_4_184 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(t_i_1_out[2])
         );
  cell_4_183 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(t_i_1_out[3])
         );
  cell_4_182 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(t_i_1_out[4])
         );
  cell_4_181 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(t_i_1_out[5])
         );
  cell_4_180 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(t_i_1_out[6])
         );
  cell_4_179 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(t_i_1_out[7])
         );
  cell_4_178 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_2_in(t_i_2_in[7]), .t_i_out(t_i_1_out[8])
         );
  cell_4_177 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[9]), .t_i_2_in(t_i_2_in[8]), .t_i_out(t_i_1_out[9])
         );
  cell_4_176 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[10]), .t_i_2_in(t_i_2_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_4_175 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[11]), .t_i_2_in(t_i_2_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_4_174 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[12]), .t_i_2_in(t_i_2_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_4_173 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[13]), .t_i_2_in(t_i_2_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_4_172 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[14]), .t_i_2_in(t_i_2_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_4_171 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[15]), .t_i_2_in(t_i_2_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_4_170 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_2_in(t_i_2_in[15]), .t_i_out(
        t_i_1_out[16]) );
  cell_4_169 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_2_in(t_i_2_in[16]), .t_i_out(
        t_i_1_out[17]) );
  cell_4_168 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_2_in(t_i_2_in[17]), .t_i_out(
        t_i_1_out[18]) );
  cell_4_167 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_2_in(t_i_2_in[18]), .t_i_out(
        t_i_1_out[19]) );
  cell_4_166 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_2_in(t_i_2_in[19]), .t_i_out(
        t_i_1_out[20]) );
  cell_4_165 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_2_in(t_i_2_in[20]), .t_i_out(
        t_i_1_out[21]) );
  cell_4_164 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_2_in(t_i_2_in[21]), .t_i_out(
        t_i_1_out[22]) );
  cell_4_163 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_2_in(t_i_2_in[22]), .t_i_out(
        t_i_1_out[23]) );
  cell_4_162 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_2_in(t_i_2_in[23]), .t_i_out(
        t_i_1_out[24]) );
  cell_4_161 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_2_in(t_i_2_in[24]), .t_i_out(
        t_i_1_out[25]) );
  cell_4_160 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_2_in(t_i_2_in[25]), .t_i_out(
        t_i_1_out[26]) );
  cell_4_159 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_2_in(t_i_2_in[26]), .t_i_out(
        t_i_1_out[27]) );
  cell_4_158 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_2_in(t_i_2_in[27]), .t_i_out(
        t_i_1_out[28]) );
  cell_4_157 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_2_in(t_i_2_in[28]), .t_i_out(
        t_i_1_out[29]) );
  cell_4_156 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_2_in(t_i_2_in[29]), .t_i_out(
        t_i_1_out[30]) );
  cell_4_155 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[31]), .t_i_2_in(t_i_2_in[30]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV2 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_185 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n1, n2;

  LVT_XOR2HSV0 U1 ( .A1(n1), .A2(n2), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n1) );
endmodule


module cell_3_5770 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5769 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5768 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5767 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5766 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5765 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5764 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5763 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5762 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5761 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5760 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5759 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5758 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5757 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5756 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5755 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5754 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5753 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5752 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5751 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5750 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5749 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5748 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5747 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5746 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5745 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5744 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5743 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5742 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5741 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV0 U2 ( .A1(n8), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2SR U3 ( .I(t_i_1_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV2 U5 ( .A1(n5), .A2(n6), .ZN(n7) );
  LVT_INHSV2 U6 ( .I(n8), .ZN(n2) );
  LVT_NAND2HSV0 U7 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XNOR2HSV4 U8 ( .A1(n9), .A2(n7), .ZN(t_i_out) );
endmodule


module cell_3_5740 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV4 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNHSV2 U4 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV0P5 U5 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2SR U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_185 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_185 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5770 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5769 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5768 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5767 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5766 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5765 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5764 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5763 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5762 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5761 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5760 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5759 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5758 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5757 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5756 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5755 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5754 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5753 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5752 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5751 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5750 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5749 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5748 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5747 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5746 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5745 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5744 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5743 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5742 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5741 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5740 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV6SR U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_184 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_5739 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5738 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5737 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5736 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5735 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5734 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5733 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5732 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5731 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5730 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5729 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5728 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5727 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5726 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5725 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5724 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5723 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5722 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5721 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5720 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5719 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5718 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5717 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5716 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5715 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5714 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
endmodule


module cell_3_5713 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_5712 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_5711 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_5710 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_CLKAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .Z(n3) );
  LVT_XNOR2HSV4 U3 ( .A1(t_i_1_in), .A2(n3), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_5709 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNHSV2P5 U1 ( .I(n7), .ZN(n4) );
  LVT_INHSV3 U2 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV8 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV4 U6 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV4 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_184 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_184 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_5739 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5738 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5737 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5736 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5735 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5734 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5733 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5732 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5731 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5730 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5729 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5728 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5727 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5726 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5725 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5724 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5723 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5722 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5721 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5720 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5719 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5718 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5717 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5716 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5715 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5714 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5713 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5712 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5711 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5710 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5709 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_183 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_5708 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5707 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5706 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5705 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5704 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5703 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5702 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5701 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5700 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5699 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5698 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5697 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5696 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5695 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5694 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5693 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5692 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5691 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5690 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5689 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5688 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5687 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5686 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5685 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5684 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5683 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5682 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5681 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5680 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5679 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_5678 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  LVT_INHSV2SR U1 ( .I(n15), .ZN(n5) );
  LVT_NAND2HSV2 U2 ( .A1(n7), .A2(n8), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U3 ( .A1(n5), .A2(n4), .ZN(n8) );
  LVT_NAND2HSV2 U4 ( .A1(n10), .A2(n13), .ZN(n11) );
  LVT_CLKNHSV2 U5 ( .I(t_i_1_in), .ZN(n10) );
  LVT_NAND2HSV2 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n15) );
  LVT_CLKNAND2HSV0 U7 ( .A1(n11), .A2(n12), .ZN(n4) );
  LVT_NAND2HSV2 U8 ( .A1(n11), .A2(n12), .ZN(n14) );
  LVT_CLKNAND2HSV0 U9 ( .A1(n9), .A2(t_i_1_in), .ZN(n12) );
  LVT_INHSV2 U10 ( .I(n14), .ZN(n6) );
  LVT_CLKNAND2HSV1 U11 ( .A1(n6), .A2(n15), .ZN(n7) );
  LVT_INHSV2 U12 ( .I(n13), .ZN(n9) );
  LVT_NAND2HSV0 U13 ( .A1(b_in), .A2(a_in), .ZN(n13) );
endmodule


module row_other_183 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_183 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_5708 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5707 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5706 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5705 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5704 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5703 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5702 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5701 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5700 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5699 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5698 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5697 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5696 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5695 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5694 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5693 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5692 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5691 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5690 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5689 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5688 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5687 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5686 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5685 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5684 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5683 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5682 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5681 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5680 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5679 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5678 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_182 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_5677 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5676 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5675 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5674 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5673 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5672 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5671 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5670 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5669 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5668 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5667 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5666 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5665 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5664 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5663 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5662 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5661 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5660 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5659 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5658 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5657 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5656 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5655 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5654 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5653 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5652 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5651 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5650 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5649 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5648 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5647 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV2 U1 ( .A1(n6), .A2(n4), .ZN(n2) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(n6), .B(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U3 ( .A1(n5), .A2(t_i_1_in), .ZN(n4) );
  LVT_CLKNAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_NAND2HSV0 U5 ( .A1(b_in), .A2(a_in), .ZN(n5) );
endmodule


module row_other_182 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_182 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5677 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5676 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5675 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5674 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5673 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5672 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5671 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5670 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5669 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5668 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5667 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5666 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5665 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5664 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5663 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5662 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5661 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5660 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5659 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5658 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5657 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5656 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5655 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5654 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5653 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5652 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5651 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5650 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5649 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5648 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5647 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2SR U1 ( .I(n2), .ZN(n3) );
  LVT_CLKNHSV0P5 U2 ( .I(t_m_1_in), .ZN(n2) );
  LVT_CLKNHSV4 U3 ( .I(n2), .ZN(n1) );
endmodule


module cell_2_181 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_5646 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5645 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5644 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5643 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5642 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5641 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5640 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5639 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5638 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5637 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5636 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5635 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5634 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5633 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5632 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5631 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5630 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5629 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5628 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5627 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5626 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5625 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5624 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5623 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5622 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5621 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5620 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5619 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5618 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5617 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_5616 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNHSV2 U2 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV3 U5 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV4 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV4 U7 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_181 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_181 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5646 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5645 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5644 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5643 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5642 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5641 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5640 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5639 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5638 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5637 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5636 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5635 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5634 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5633 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5632 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5631 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5630 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5629 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5628 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5627 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5626 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5625 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5624 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5623 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5622 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5621 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5620 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5619 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5618 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5617 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5616 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_180 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_5615 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5614 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5613 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5612 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5611 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5610 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5609 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5608 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5607 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5606 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5605 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5604 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5603 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5602 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5601 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5600 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5599 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5598 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5597 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5596 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5595 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5594 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5593 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5592 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5591 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5590 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5589 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5588 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV0 U4 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV1 U5 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_5587 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5586 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5585 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U1 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_INHSV2SR U2 ( .I(n10), .ZN(n4) );
  LVT_XOR2HSV2 U4 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_NAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_CLKNHSV0P5 U6 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV0P5 U7 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_NAND2HSV2 U8 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
endmodule


module row_other_180 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_180 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5615 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5614 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5613 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5612 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5611 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5610 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5609 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5608 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5607 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5606 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5605 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5604 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5603 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5602 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5601 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5600 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5599 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5598 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5597 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5596 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5595 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5594 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5593 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5592 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5591 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5590 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5589 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5588 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5587 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5586 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5585 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n3) );
  LVT_INHSV2 U2 ( .I(n3), .ZN(n1) );
  LVT_INHSV2 U3 ( .I(n3), .ZN(n2) );
endmodule


module cell_2_179 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_5584 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5583 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5582 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5581 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5580 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5579 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5578 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5577 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5576 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5575 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5574 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5573 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5572 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5571 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5570 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5569 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5568 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5567 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5566 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5565 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5564 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5563 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5562 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5561 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5560 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5559 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5558 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5557 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5556 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5555 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5554 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_NAND2HSV3 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV2 U2 ( .I(n9), .ZN(n4) );
  LVT_CLKNAND2HSV1 U3 ( .A1(n4), .A2(n2), .ZN(n6) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XOR2HSV0 U5 ( .A1(n8), .A2(t_i_1_in), .Z(n2) );
  LVT_NAND2HSV0 U6 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U7 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_XNOR2HSV1 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_179 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_2_179 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5584 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5583 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5582 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5581 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5580 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5579 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5578 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5577 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5576 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5575 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5574 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5573 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5572 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5571 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5570 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5569 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5568 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5567 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5566 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5565 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5564 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5563 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5562 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5561 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5560 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5559 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5558 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5557 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5556 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5555 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5554 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV1 U1 ( .I(n3), .ZN(n4) );
  LVT_INHSV0P5SR U2 ( .I(t_m_1_in), .ZN(n3) );
  LVT_INHSV0SR U3 ( .I(n3), .ZN(n1) );
  LVT_INHSV0SR U4 ( .I(n3), .ZN(n2) );
endmodule


module cell_2_178 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_5553 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5552 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5551 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5550 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5549 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5548 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5547 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5546 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5545 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5544 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5543 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5542 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5541 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5540 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5539 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5538 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5537 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5536 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5535 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5534 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5533 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5532 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5531 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5530 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5529 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5528 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5527 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_5526 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5525 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5524 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5523 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV1 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_178 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_178 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_5553 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5552 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5551 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5550 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5549 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5548 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5547 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5546 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5545 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5544 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5543 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5542 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5541 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5540 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5539 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5538 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5537 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5536 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5535 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5534 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5533 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5532 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5531 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5530 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5529 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5528 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5527 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5526 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5525 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5524 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5523 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_CLKNHSV0P5 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_177 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_5522 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5521 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5520 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5519 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5518 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5517 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5516 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5515 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5514 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5513 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5512 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5511 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5510 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5509 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5508 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5507 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5506 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5505 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5504 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5503 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5502 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5501 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5500 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5499 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5498 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5497 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5496 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV3 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5495 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5494 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5493 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_5492 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_IOA21HSV4 U1 ( .A1(n8), .A2(n6), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV3 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKNHSV2P5 U4 ( .I(n6), .ZN(n4) );
  LVT_XNOR2HSV4 U5 ( .A1(n7), .A2(t_i_1_in), .ZN(n6) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n2), .A2(n4), .ZN(n5) );
  LVT_INHSV2 U7 ( .I(n8), .ZN(n2) );
endmodule


module row_other_177 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_2_177 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5522 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5521 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5520 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5519 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5518 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5517 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5516 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5515 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5514 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5513 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5512 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5511 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5510 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5509 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5508 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5507 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5506 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5505 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5504 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5503 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5502 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5501 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5500 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5499 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5498 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5497 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5496 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5495 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5494 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5493 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5492 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV6 U1 ( .I(n4), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n3), .ZN(n4) );
  LVT_INHSV2 U3 ( .I(t_m_1_in), .ZN(n2) );
  LVT_INHSV4SR U4 ( .I(n2), .ZN(n3) );
endmodule


module cell_2_176 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_5491 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5490 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5489 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5488 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5487 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5486 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5485 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5484 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5483 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5482 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5481 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5480 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5479 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5478 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5477 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5476 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5475 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5474 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5473 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5472 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5471 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5470 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5469 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5468 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5467 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5466 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5465 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5464 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_5463 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5462 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5461 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2SR U2 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV2 U4 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNAND2HSV0 U5 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV3 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV4 U7 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_INHSV2 U8 ( .I(n7), .ZN(n4) );
endmodule


module row_other_176 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_176 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5491 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5490 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5489 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5488 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5487 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5486 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5485 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5484 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5483 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5482 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5481 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5480 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5479 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5478 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5477 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5476 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5475 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5474 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5473 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5472 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5471 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5470 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5469 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5468 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5467 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5466 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5465 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5464 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5463 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5462 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5461 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV4 U1 ( .I(n2), .ZN(n1) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n2) );
endmodule


module cell_2_175 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_5460 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5459 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5458 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5457 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5456 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5455 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5454 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5453 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5452 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5451 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5450 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5449 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5448 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5447 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5446 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5445 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5444 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5443 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5442 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5441 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5440 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5439 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5438 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5437 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U4 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U5 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_5436 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5435 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5434 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5433 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5432 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5431 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5430 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV4 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV4SR U4 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV3 U5 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U6 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
  LVT_NAND2HSV4 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV2 U8 ( .I(n7), .ZN(n4) );
endmodule


module row_other_175 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_175 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5460 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5459 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5458 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5457 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5456 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5455 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5454 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5453 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5452 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5451 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5450 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5449 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5448 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5447 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5446 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5445 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5444 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5443 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5442 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5441 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5440 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5439 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5438 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5437 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5436 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5435 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5434 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5433 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5432 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5431 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5430 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_174 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_5429 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5428 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5427 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5426 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5425 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5424 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5423 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5422 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5421 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5420 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5419 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5418 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5417 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5416 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5415 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5414 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5413 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5412 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5411 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5410 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5409 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5408 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5407 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5406 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5405 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5404 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_5403 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5402 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5401 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5400 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5399 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_CLKNHSV2 U2 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_CLKNHSV2 U5 ( .I(n10), .ZN(n4) );
  LVT_XOR2HSV2 U6 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_NAND2HSV2 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_CLKNAND2HSV1 U8 ( .A1(n10), .A2(n5), .ZN(n6) );
endmodule


module row_other_174 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_2_174 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5429 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5428 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5427 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5426 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5425 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5424 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5423 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5422 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5421 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5420 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5419 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5418 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5417 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5416 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5415 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5414 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5413 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5412 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5411 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5410 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5409 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5408 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5407 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5406 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5405 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5404 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5403 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5402 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5401 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5400 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5399 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV4SR U1 ( .I(n1), .ZN(n3) );
  LVT_INHSV4SR U2 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV0P5SR U3 ( .I(n1), .ZN(n2) );
  LVT_INHSV2P5 U4 ( .I(n1), .ZN(n4) );
endmodule


module cell_2_173 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_5398 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5397 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5396 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5395 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5394 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5393 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5392 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5391 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5390 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5389 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5388 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5387 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5386 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5385 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5384 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5383 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5382 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5381 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5380 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5379 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5378 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5377 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5376 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5375 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5374 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5373 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5372 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5371 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5370 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5369 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_CLKNHSV0P5 U5 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_5368 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9, n10;

  LVT_OAI21HSV2 U1 ( .A1(t_i_1_in), .A2(n9), .B(n2), .ZN(n8) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_CLKNAND2HSV0 U3 ( .A1(n9), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n9) );
  LVT_NAND2HSV0 U5 ( .A1(n10), .A2(n8), .ZN(n6) );
  LVT_NAND2HSV2 U6 ( .A1(n7), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U7 ( .A1(n4), .A2(n5), .ZN(n7) );
  LVT_INHSV2SR U8 ( .I(n10), .ZN(n4) );
  LVT_INHSV2 U9 ( .I(n8), .ZN(n5) );
endmodule


module row_other_173 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_173 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5398 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5397 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5396 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5395 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5394 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5393 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5392 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5391 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5390 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5389 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5388 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5387 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5386 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5385 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5384 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5383 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5382 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5381 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5380 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5379 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5378 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5377 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5376 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5375 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5374 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5373 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5372 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5371 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5370 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5369 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5368 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV6 U1 ( .I(n2), .ZN(n3) );
  LVT_INHSV2SR U2 ( .I(t_m_1_in), .ZN(n2) );
  LVT_CLKNHSV2 U3 ( .I(n2), .ZN(n1) );
endmodule


module cell_2_172 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_5367 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5366 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5365 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5364 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5363 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5362 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5361 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5360 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5359 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5358 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5357 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5356 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5355 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5354 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5353 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5352 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5351 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5350 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5349 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5348 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5347 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5346 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5345 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5344 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5343 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5342 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_5341 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_5340 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5339 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n5), .A2(n6), .Z(t_i_out) );
endmodule


module cell_3_5338 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_5337 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_OAI21HSV2 U2 ( .A1(n2), .A2(n6), .B(n4), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U3 ( .A1(t_i_1_in), .A2(n5), .ZN(n2) );
  LVT_CLKNAND2HSV1 U4 ( .A1(n2), .A2(n6), .ZN(n4) );
  LVT_NAND2HSV0 U5 ( .A1(b_in), .A2(a_in), .ZN(n5) );
endmodule


module row_other_172 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_172 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5367 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5366 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5365 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5364 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5363 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5362 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5361 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5360 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5359 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5358 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5357 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5356 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5355 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5354 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5353 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5352 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5351 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5350 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5349 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5348 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5347 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5346 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5345 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5344 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5343 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5342 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5341 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5340 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5339 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5338 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5337 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV6SR U1 ( .I(n2), .ZN(n3) );
  LVT_CLKNHSV2 U2 ( .I(t_m_1_in), .ZN(n2) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
endmodule


module cell_2_171 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_5336 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5335 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5334 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5333 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5332 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5331 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5330 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5329 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5328 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5327 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5326 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5325 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5324 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5323 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5322 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5321 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5320 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5319 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5318 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5317 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5316 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5315 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5314 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5313 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5312 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5311 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_5310 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_5309 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5308 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5307 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5306 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_171 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_171 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5336 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5335 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5334 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5333 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5332 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5331 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5330 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5329 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5328 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5327 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5326 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5325 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5324 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5323 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5322 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5321 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5320 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5319 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5318 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5317 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5316 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5315 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5314 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5313 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5312 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5311 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5310 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5309 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5308 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5307 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5306 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV10SR U1 ( .I(n3), .ZN(n2) );
  LVT_CLKNHSV6 U2 ( .I(t_m_1_in), .ZN(n3) );
  LVT_INHSV2 U3 ( .I(n3), .ZN(n1) );
endmodule


module cell_2_170 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_5305 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5304 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5303 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5302 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5301 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5300 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5299 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5298 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5297 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5296 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5295 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5294 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5293 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5292 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5291 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5290 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5289 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5288 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5287 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5286 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5285 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5284 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5283 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5282 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5281 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5280 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5279 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5278 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_5277 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5276 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5275 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_CLKNAND2HSV2 U1 ( .A1(n6), .A2(n4), .ZN(n2) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(t_i_1_in), .ZN(n4) );
  LVT_OAI21HSV2 U4 ( .A1(n6), .A2(n4), .B(n2), .ZN(t_i_out) );
  LVT_CLKNAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module row_other_170 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_170 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_5305 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5304 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5303 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5302 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5301 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5300 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5299 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5298 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5297 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5296 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5295 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5294 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5293 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5292 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5291 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5290 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5289 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5288 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5287 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5286 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5285 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5284 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5283 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5282 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5281 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5280 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5279 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5278 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5277 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5276 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5275 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_169 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_5274 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5273 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5272 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5271 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5270 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5269 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5268 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5267 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5266 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5265 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5264 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5263 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5262 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5261 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5260 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5259 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5258 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5257 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5256 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5255 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5254 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5253 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5252 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5251 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5250 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5249 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5248 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5247 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5246 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5245 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5244 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV2 U2 ( .I(n9), .ZN(n2) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
  LVT_NAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV0P5 U7 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2 U8 ( .I(n7), .ZN(n4) );
endmodule


module row_other_169 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_169 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5274 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5273 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5272 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5271 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5270 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5269 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5268 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5267 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5266 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5265 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5264 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5263 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5262 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5261 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5260 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5259 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5258 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5257 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5256 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5255 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5254 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5253 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5252 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5251 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5250 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5249 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5248 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5247 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5246 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5245 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5244 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV6 U1 ( .I(n2), .ZN(n3) );
  LVT_CLKNHSV2 U2 ( .I(t_m_1_in), .ZN(n2) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
endmodule


module cell_2_168 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_5243 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5242 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5241 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5240 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5239 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5238 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5237 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5236 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5235 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5234 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5233 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5232 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5231 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5230 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5229 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5228 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5227 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5226 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5225 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5224 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5223 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5222 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5221 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5220 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5219 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_5218 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5217 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5216 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5215 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV2 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0P5 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNAND2HSV3 U3 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_CLKNHSV0 U4 ( .I(n8), .ZN(n4) );
  LVT_CLKNHSV2 U5 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV0 U6 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_XOR2HSV4 U8 ( .A1(n10), .A2(n9), .Z(t_i_out) );
endmodule


module cell_3_5214 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_5213 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module row_other_168 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_168 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5243 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5242 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5241 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5240 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5239 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5238 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5237 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5236 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5235 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5234 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5233 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5232 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5231 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5230 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5229 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5228 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5227 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5226 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5225 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5224 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5223 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5222 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5221 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5220 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5219 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5218 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5217 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5216 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5215 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5214 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5213 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV5 U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_CLKNHSV12 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_167 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_5212 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5211 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5210 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5209 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5208 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5207 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5206 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5205 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5204 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5203 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5202 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5201 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5200 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5199 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5198 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5197 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5196 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5195 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5194 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5193 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5192 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5191 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5190 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5189 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5188 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5187 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5186 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5185 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5184 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5183 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_CLKAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .Z(n3) );
  LVT_XNOR2HSV4 U4 ( .A1(n3), .A2(t_i_1_in), .ZN(n4) );
endmodule


module cell_3_5182 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV0 U2 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV2 U4 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV2 U5 ( .I(n9), .ZN(n2) );
  LVT_INHSV2SR U6 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV2 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_167 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_167 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5212 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5211 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5210 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5209 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5208 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5207 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5206 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5205 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5204 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5203 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5202 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5201 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5200 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5199 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5198 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5197 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5196 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5195 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5194 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5193 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5192 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5191 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5190 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5189 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5188 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5187 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5186 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5185 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5184 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5183 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5182 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2P5 U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV12SR U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_166 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_5181 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5180 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5179 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5178 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5177 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5176 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5175 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5174 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5173 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5172 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5171 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5170 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5169 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5168 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5167 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5166 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5165 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5164 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5163 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5162 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5161 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5160 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5159 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5158 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5157 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5156 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5155 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5154 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_5153 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5152 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5151 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_INAND2HSV0 U1 ( .A1(n8), .B1(n9), .ZN(n5) );
  LVT_INHSV3SR U2 ( .I(n9), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XOR2HSV0 U6 ( .A1(n7), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV2 U7 ( .A1(n4), .A2(n8), .ZN(n6) );
endmodule


module row_other_166 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_166 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5181 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5180 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5179 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5178 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5177 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5176 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5175 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5174 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5173 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5172 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5171 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5170 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5169 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5168 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5167 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5166 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5165 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5164 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5163 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5162 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5161 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5160 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5159 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5158 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5157 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5156 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5155 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5154 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5153 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5152 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5151 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV6 U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV12SR U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_165 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_5150 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5149 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5148 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5147 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5146 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5145 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5144 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5143 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5142 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5141 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5140 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5139 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5138 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5137 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5136 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5135 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5134 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5133 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5132 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5131 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5130 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5129 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5128 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5127 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5126 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5125 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5124 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5123 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5122 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5121 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_NAND2HSV0P5 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_CLKNHSV0P5 U4 ( .I(n10), .ZN(n4) );
  LVT_NAND2HSV0P5 U5 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U6 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_CLKNHSV2 U7 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV0 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_5120 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module row_other_165 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_165 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_5150 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5149 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5148 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5147 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5146 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5145 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5144 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5143 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5142 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5141 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5140 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5139 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5138 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5137 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5136 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5135 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5134 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5133 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5132 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5131 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5130 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5129 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5128 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5127 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5126 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5125 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5124 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5123 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5122 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5121 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5120 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_164 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_5119 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5118 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5117 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5116 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5115 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5114 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5113 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5112 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5111 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5110 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5109 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5108 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5107 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5106 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5105 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5104 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5103 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5102 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5101 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5100 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5099 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5098 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5097 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5096 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5095 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5094 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5093 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_5092 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_5091 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5090 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_5089 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U2 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV1 U5 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV0P5 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2 U7 ( .I(n9), .ZN(n2) );
  LVT_INHSV2 U8 ( .I(n7), .ZN(n4) );
endmodule


module row_other_164 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_164 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5119 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5118 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5117 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5116 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5115 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5114 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5113 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5112 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5111 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5110 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5109 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5108 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5107 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5106 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5105 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5104 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5103 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5102 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5101 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5100 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5099 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5098 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5097 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5096 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5095 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5094 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5093 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5092 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5091 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5090 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5089 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2 U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV12SR U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_163 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_5088 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5087 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5086 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5085 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5084 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5083 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5082 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5081 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5080 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5079 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5078 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5077 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5076 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5075 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5074 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5073 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5072 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5071 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5070 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5069 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5068 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5067 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5066 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5065 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5064 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5063 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5062 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_5061 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5060 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5059 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5058 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module row_other_163 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_163 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5088 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5087 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5086 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5085 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5084 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5083 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5082 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5081 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5080 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5079 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5078 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5077 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5076 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5075 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5074 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5073 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5072 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5071 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5070 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5069 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5068 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5067 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5066 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5065 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5064 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5063 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5062 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5061 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5060 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5059 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5058 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV6 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV4SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_162 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_5057 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5056 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5055 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5054 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5053 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5052 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5051 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5050 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5049 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5048 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5047 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5046 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5045 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5044 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5043 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5042 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5041 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5040 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5039 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5038 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5037 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5036 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5035 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5034 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5033 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5032 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5031 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5030 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5029 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5028 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5027 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV2SR U1 ( .I(n9), .ZN(n2) );
  LVT_XNOR2HSV1 U2 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_INHSV2 U4 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV1 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV4 U8 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
endmodule


module row_other_162 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_2_162 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5057 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5056 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5055 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5054 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5053 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5052 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5051 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5050 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5049 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5048 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5047 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5046 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5045 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5044 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5043 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5042 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5041 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5040 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5039 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5038 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5037 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5036 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5035 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5034 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5033 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5032 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5031 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_5030 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_5029 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_5028 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_5027 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2 U1 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U2 ( .I(n3), .ZN(n1) );
  LVT_CLKNHSV2 U3 ( .I(t_m_1_in), .ZN(n3) );
  LVT_INHSV0P5SR U4 ( .I(n3), .ZN(n4) );
endmodule


module cell_2_161 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_5026 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5025 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5024 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5023 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5022 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5021 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_5020 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_5019 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5018 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5017 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5016 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5015 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5014 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5013 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5012 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5011 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5010 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5009 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5008 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5007 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5006 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5005 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5004 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5003 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5002 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5001 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_5000 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4999 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4998 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4997 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4996 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2SR U2 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV2 U4 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U5 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U6 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
  LVT_INHSV2 U7 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV1 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
endmodule


module row_other_161 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_161 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_5026 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_5025 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_5024 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_5023 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_5022 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_5021 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_5020 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_5019 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_5018 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_5017 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_5016 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_5015 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_5014 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_5013 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_5012 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_5011 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_5010 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_5009 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_5008 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_5007 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_5006 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_5005 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_5004 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_5003 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_5002 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5001 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_5000 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4999 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4998 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4997 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4996 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV3 U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_CLKNHSV12 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_160 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_4995 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4994 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4993 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4992 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4991 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4990 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4989 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4988 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4987 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4986 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4985 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4984 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4983 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4982 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4981 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4980 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4979 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4978 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4977 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4976 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4975 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4974 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4973 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4972 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4971 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4970 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4969 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4968 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4967 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4966 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4965 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n2), .A2(n4), .ZN(n5) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNHSV2 U4 ( .I(n9), .ZN(n2) );
  LVT_CLKNHSV3 U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV1 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV1 U7 ( .A1(n9), .A2(n7), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_160 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_160 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4995 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4994 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4993 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4992 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4991 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4990 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4989 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4988 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4987 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4986 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4985 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4984 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4983 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4982 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4981 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4980 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4979 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4978 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4977 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4976 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4975 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4974 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4973 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4972 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4971 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4970 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4969 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4968 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4967 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4966 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4965 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV3 U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_CLKNHSV12 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_159 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_4964 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4963 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4962 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4961 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4960 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4959 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4958 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4957 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4956 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4955 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4954 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4953 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4952 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4951 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4950 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4949 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4948 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4947 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4946 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4945 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4944 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4943 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4942 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4941 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4940 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4939 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4938 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4937 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV0P5 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_4936 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4935 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_XOR2HSV0 U2 ( .A1(n7), .A2(n8), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U3 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV0 U5 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_3_4934 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_IOA21HSV4 U1 ( .A1(n2), .A2(n4), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(n8), .A2(n6), .ZN(n5) );
  LVT_CLKNHSV2 U4 ( .I(n8), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n6), .ZN(n4) );
  LVT_CLKNAND2HSV1 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XNOR2HSV1 U7 ( .A1(t_i_1_in), .A2(n7), .ZN(n6) );
endmodule


module row_other_159 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_159 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4964 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4963 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4962 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4961 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4960 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4959 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4958 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4957 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4956 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4955 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4954 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4953 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4952 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4951 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4950 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4949 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4948 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4947 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4946 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4945 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4944 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4943 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4942 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4941 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4940 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4939 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4938 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4937 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4936 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4935 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4934 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV8 U1 ( .I(n2), .ZN(n1) );
  LVT_INHSV2P5 U2 ( .I(t_m_1_in), .ZN(n2) );
endmodule


module cell_2_158 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4933 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4932 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4931 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4930 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4929 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4928 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4927 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4926 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4925 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4924 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4923 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4922 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4921 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4920 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4919 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4918 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4917 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4916 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4915 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4914 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4913 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4912 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4911 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4910 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4909 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4908 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4907 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4906 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4905 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4904 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4903 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_158 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_2_158 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_4933 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4932 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4931 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4930 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4929 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4928 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4927 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4926 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4925 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4924 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4923 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4922 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4921 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4920 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4919 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4918 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4917 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4916 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4915 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4914 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4913 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4912 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4911 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4910 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4909 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4908 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4907 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4906 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4905 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4904 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4903 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV8 U1 ( .I(t_m_1_in), .Z(n1) );
  LVT_CLKBUFHSV4 U2 ( .I(t_m_1_in), .Z(n2) );
  LVT_INHSV0SR U3 ( .I(t_m_1_in), .ZN(n3) );
  LVT_INHSV0P5SR U4 ( .I(n3), .ZN(n4) );
endmodule


module cell_2_157 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4902 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4901 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4900 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4899 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4898 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4897 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4896 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4895 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4894 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4893 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4892 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4891 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4890 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4889 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4888 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4887 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4886 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4885 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4884 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4883 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4882 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4881 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4880 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4879 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4878 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4877 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4876 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4875 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4874 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4873 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4872 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2P5 U5 ( .I(n9), .ZN(n2) );
  LVT_INHSV3 U6 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV2 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_157 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_157 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_4902 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4901 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4900 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4899 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4898 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4897 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4896 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4895 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4894 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4893 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4892 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4891 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4890 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4889 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4888 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4887 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4886 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4885 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4884 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4883 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4882 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4881 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4880 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4879 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4878 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4877 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4876 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4875 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4874 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4873 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4872 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV4SR U1 ( .I(t_m_1_in), .ZN(n2) );
  LVT_CLKNHSV8 U2 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n3) );
endmodule


module cell_2_156 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_4871 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4870 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4869 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4868 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4867 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4866 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4865 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4864 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4863 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4862 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4861 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4860 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4859 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4858 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4857 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4856 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4855 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4854 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4853 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4852 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4851 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4850 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4849 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4848 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4847 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4846 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4845 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4844 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4843 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4842 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4841 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_156 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_156 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_4871 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4870 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4869 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4868 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4867 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4866 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4865 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4864 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4863 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4862 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4861 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4860 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4859 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4858 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4857 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4856 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4855 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4854 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4853 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4852 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4851 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4850 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4849 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4848 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4847 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4846 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4845 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4844 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4843 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4842 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4841 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_155 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_4840 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4839 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4838 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4837 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV1 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_4836 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4835 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4834 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4833 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4832 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4831 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_4830 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4829 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4828 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4827 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_4826 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4825 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4824 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4823 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4822 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4821 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4820 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4819 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4818 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4817 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4816 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4815 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4814 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4813 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4812 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4811 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV1 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_4810 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(t_i_1_in), .ZN(n4) );
  LVT_OAI21HSV0 U2 ( .A1(n6), .A2(n4), .B(n2), .ZN(t_i_out) );
  LVT_CLKNAND2HSV0 U5 ( .A1(n6), .A2(n4), .ZN(n2) );
endmodule


module row_other_155 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_155 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_4840 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4839 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4838 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4837 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4836 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4835 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4834 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4833 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4832 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4831 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4830 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4829 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4828 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4827 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4826 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4825 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4824 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4823 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4822 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4821 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4820 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4819 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4818 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4817 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4816 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4815 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4814 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4813 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4812 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4811 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4810 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_5 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [31:0] a_in;
  input [31:0] g_in;
  input [31:0] b_in;
  input [31:0] t_m_1_in;
  input [30:0] t_i_1_in;
  input [30:0] t_i_2_in;
  output [31:0] a_out;
  output [31:0] g_out;
  output [30:0] t_i_1_out;
  output [30:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;
  wire   n1, n2, n4, n5, n7, n8, n10, n11, n12, n13, n14;
  wire   [30:0] t0;
  wire   [30:0] t1;
  wire   [30:0] t2;
  wire   [30:0] t3;
  wire   [30:0] t4;
  wire   [30:0] t5;
  wire   [30:0] t6;
  wire   [30:0] t7;
  wire   [30:0] t8;
  wire   [30:0] t9;
  wire   [30:0] t10;
  wire   [30:0] t11;
  wire   [30:0] t12;
  wire   [30:0] t13;
  wire   [30:0] t14;
  wire   [30:0] t15;
  wire   [30:0] t16;
  wire   [30:0] t17;
  wire   [30:0] t18;
  wire   [30:0] t19;
  wire   [30:0] t20;
  wire   [30:0] t21;
  wire   [30:0] t22;
  wire   [30:0] t23;
  wire   [30:0] t24;
  wire   [30:0] t25;
  wire   [30:0] t26;
  wire   [30:0] t27;
  wire   [30:0] t28;
  wire   [30:0] t29;
  wire   [30:0] t30;
  assign a_out[31] = a_in[31];
  assign a_out[30] = a_in[30];
  assign a_out[29] = a_in[29];
  assign a_out[28] = a_in[28];
  assign a_out[27] = a_in[27];
  assign a_out[26] = a_in[26];
  assign a_out[25] = a_in[25];
  assign a_out[24] = a_in[24];
  assign a_out[22] = a_in[22];
  assign a_out[21] = a_in[21];
  assign a_out[18] = a_in[18];
  assign a_out[17] = a_in[17];
  assign a_out[16] = a_in[16];
  assign a_out[15] = a_in[15];
  assign a_out[14] = a_in[14];
  assign a_out[13] = a_in[13];
  assign a_out[12] = a_in[12];
  assign a_out[11] = a_in[11];
  assign a_out[10] = a_in[10];
  assign a_out[9] = a_in[9];
  assign a_out[8] = a_in[8];
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[30] = g_in[30];
  assign g_out[29] = g_in[29];
  assign g_out[28] = g_in[28];
  assign g_out[27] = g_in[27];
  assign g_out[26] = g_in[26];
  assign g_out[25] = g_in[25];
  assign g_out[24] = g_in[24];
  assign g_out[23] = g_in[23];
  assign g_out[22] = g_in[22];
  assign g_out[21] = g_in[21];
  assign g_out[20] = g_in[20];
  assign g_out[19] = g_in[19];
  assign g_out[18] = g_in[18];
  assign g_out[17] = g_in[17];
  assign g_out[16] = g_in[16];
  assign g_out[15] = g_in[15];
  assign g_out[14] = g_in[14];
  assign g_out[13] = g_in[13];
  assign g_out[12] = g_in[12];
  assign g_out[11] = g_in[11];
  assign g_out[10] = g_in[10];
  assign g_out[9] = g_in[9];
  assign g_out[8] = g_in[8];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_5 u0 ( .a_in({a_in[31:24], n5, a_in[22:21], n2, n8, a_in[18:0]}), 
        .g_in(g_in), .b_in(b_in[31]), .t_m_1_in(t_m_1_in[31]), .t_i_1_in({
        t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), .t_i_1_out(t0), 
        .t_i_2_out(t_i_2_out[30]) );
  row_other_185 u1 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in(g_in), .b_in(b_in[30]), .t_m_1_in(t_m_1_in[30]), 
        .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[29]) );
  row_other_184 u2 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in(g_in), .b_in(b_in[29]), .t_m_1_in(t_m_1_in[29]), 
        .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[28]) );
  row_other_183 u3 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in(g_in), .b_in(b_in[28]), .t_m_1_in(t_m_1_in[28]), 
        .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[27]) );
  row_other_182 u4 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[27]), 
        .t_m_1_in(t_m_1_in[27]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(
        t_i_2_out[26]) );
  row_other_181 u5 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[26]), 
        .t_m_1_in(n13), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(
        t_i_2_out[25]) );
  row_other_180 u6 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[25]), 
        .t_m_1_in(t_m_1_in[25]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(
        t_i_2_out[24]) );
  row_other_179 u7 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[24]), 
        .t_m_1_in(t_m_1_in[24]), .t_i_1_in(t6), .t_i_1_out(t7), .t_i_2_out(
        t_i_2_out[23]) );
  row_other_178 u8 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[23]), 
        .t_m_1_in(t_m_1_in[23]), .t_i_1_in(t7), .t_i_1_out(t8), .t_i_2_out(
        t_i_2_out[22]) );
  row_other_177 u9 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[22]), 
        .t_m_1_in(t_m_1_in[22]), .t_i_1_in(t8), .t_i_1_out(t9), .t_i_2_out(
        t_i_2_out[21]) );
  row_other_176 u10 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[21]), 
        .t_m_1_in(t_m_1_in[21]), .t_i_1_in(t9), .t_i_1_out(t10), .t_i_2_out(
        t_i_2_out[20]) );
  row_other_175 u11 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[20]), 
        .t_m_1_in(t_m_1_in[20]), .t_i_1_in(t10), .t_i_1_out(t11), .t_i_2_out(
        t_i_2_out[19]) );
  row_other_174 u12 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[19]), 
        .t_m_1_in(t_m_1_in[19]), .t_i_1_in(t11), .t_i_1_out(t12), .t_i_2_out(
        t_i_2_out[18]) );
  row_other_173 u13 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[18]), 
        .t_m_1_in(t_m_1_in[18]), .t_i_1_in(t12), .t_i_1_out(t13), .t_i_2_out(
        t_i_2_out[17]) );
  row_other_172 u14 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[17]), 
        .t_m_1_in(t_m_1_in[17]), .t_i_1_in(t13), .t_i_1_out(t14), .t_i_2_out(
        t_i_2_out[16]) );
  row_other_171 u15 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[16]), 
        .t_m_1_in(t_m_1_in[16]), .t_i_1_in(t14), .t_i_1_out(t15), .t_i_2_out(
        t_i_2_out[15]) );
  row_other_170 u16 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[15]), 
        .t_m_1_in(n11), .t_i_1_in(t15), .t_i_1_out(t16), .t_i_2_out(
        t_i_2_out[14]) );
  row_other_169 u17 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[14]), 
        .t_m_1_in(t_m_1_in[14]), .t_i_1_in(t16), .t_i_1_out(t17), .t_i_2_out(
        t_i_2_out[13]) );
  row_other_168 u18 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[13]), 
        .t_m_1_in(t_m_1_in[13]), .t_i_1_in(t17), .t_i_1_out(t18), .t_i_2_out(
        t_i_2_out[12]) );
  row_other_167 u19 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[12]), 
        .t_m_1_in(t_m_1_in[12]), .t_i_1_in(t18), .t_i_1_out(t19), .t_i_2_out(
        t_i_2_out[11]) );
  row_other_166 u20 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[11]), 
        .t_m_1_in(t_m_1_in[11]), .t_i_1_in(t19), .t_i_1_out(t20), .t_i_2_out(
        t_i_2_out[10]) );
  row_other_165 u21 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[10]), 
        .t_m_1_in(t_m_1_in[10]), .t_i_1_in(t20), .t_i_1_out(t21), .t_i_2_out(
        t_i_2_out[9]) );
  row_other_164 u22 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[9]), 
        .t_m_1_in(t_m_1_in[9]), .t_i_1_in(t21), .t_i_1_out(t22), .t_i_2_out(
        t_i_2_out[8]) );
  row_other_163 u23 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[8]), 
        .t_m_1_in(t_m_1_in[8]), .t_i_1_in(t22), .t_i_1_out(t23), .t_i_2_out(
        t_i_2_out[7]) );
  row_other_162 u24 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[7]), 
        .t_m_1_in(t_m_1_in[7]), .t_i_1_in(t23), .t_i_1_out(t24), .t_i_2_out(
        t_i_2_out[6]) );
  row_other_161 u25 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[6]), 
        .t_m_1_in(t_m_1_in[6]), .t_i_1_in(t24), .t_i_1_out(t25), .t_i_2_out(
        t_i_2_out[5]) );
  row_other_160 u26 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[5]), 
        .t_m_1_in(t_m_1_in[5]), .t_i_1_in(t25), .t_i_1_out(t26), .t_i_2_out(
        t_i_2_out[4]) );
  row_other_159 u27 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[4]), 
        .t_m_1_in(t_m_1_in[4]), .t_i_1_in(t26), .t_i_1_out(t27), .t_i_2_out(
        t_i_2_out[3]) );
  row_other_158 u28 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[3]), 
        .t_m_1_in(t_m_1_in[3]), .t_i_1_in(t27), .t_i_1_out(t28), .t_i_2_out(
        t_i_2_out[2]) );
  row_other_157 u29 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[2]), 
        .t_m_1_in(t_m_1_in[2]), .t_i_1_in(t28), .t_i_1_out(t29), .t_i_2_out(
        t_i_2_out[1]) );
  row_other_156 u30 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[1]), 
        .t_m_1_in(t_m_1_in[1]), .t_i_1_in(t29), .t_i_1_out(t30), .t_i_2_out(
        t_i_2_out[0]) );
  row_other_155 u31 ( .a_in({a_in[31:24], a_out[23], a_in[22:21], a_out[20:19], 
        a_in[18:0]}), .g_in({g_out[31], g_in[30:0]}), .b_in(b_in[0]), 
        .t_m_1_in(t_m_1_in[0]), .t_i_1_in(t30), .t_i_1_out(t_i_1_out), 
        .t_i_2_out(t_i_1_out_0) );
  LVT_INHSV2 U1 ( .I(a_in[19]), .ZN(n7) );
  LVT_INHSV2 U2 ( .I(a_in[20]), .ZN(n1) );
  LVT_INHSV2 U3 ( .I(a_in[23]), .ZN(n4) );
  LVT_CLKNHSV8 U4 ( .I(t_m_1_in[15]), .ZN(n10) );
  LVT_INHSV2SR U5 ( .I(n1), .ZN(n2) );
  LVT_INHSV2SR U6 ( .I(n1), .ZN(a_out[20]) );
  LVT_INHSV2SR U7 ( .I(n4), .ZN(n5) );
  LVT_INHSV2SR U8 ( .I(n4), .ZN(a_out[23]) );
  LVT_CLKNHSV2 U9 ( .I(n7), .ZN(n8) );
  LVT_INHSV2SR U10 ( .I(n7), .ZN(a_out[19]) );
  LVT_INHSV10 U11 ( .I(n12), .ZN(n13) );
  LVT_INHSV4 U12 ( .I(t_m_1_in[26]), .ZN(n12) );
  LVT_CLKNHSV4 U13 ( .I(n14), .ZN(g_out[31]) );
  LVT_INHSV12SR U14 ( .I(n10), .ZN(n11) );
  LVT_INHSV0SR U15 ( .I(g_in[31]), .ZN(n14) );
endmodule


module regist_32bit_31 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_32bit_30 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_31bit_20 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n2), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n2), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n2), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n1), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module PE_5 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro );
  input [31:0] a_in;
  input [31:0] g_in;
  input [31:0] b_in;
  input [30:0] t_i_1_in;
  input [30:0] t_i_2_in;
  output [31:0] a_out;
  output [31:0] g_out;
  output [31:0] b_out;
  output [30:0] t_i_1_out;
  output [30:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   n80, l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n71, n72, n73,
         n74, n75, n76, n77, n78, n79;
  wire   [31:0] l_a;
  wire   [31:0] l_g;
  wire   [30:0] l_t_i_1_in;
  wire   [30:0] l_t_i_2_in;
  wire   [31:0] mux_b;
  wire   [31:0] mux_bq;
  wire   [30:0] to_7;
  wire   [30:0] ti_7;
  wire   [31:0] ao;
  wire   [31:0] go;
  wire   [30:0] to;

  LVT_AO22HSV0 U35 ( .A1(mux_bq[9]), .A2(n35), .B1(b_out[9]), .B2(n26), .Z(
        mux_b[9]) );
  LVT_AO22HSV0 U36 ( .A1(mux_bq[8]), .A2(n35), .B1(b_out[8]), .B2(n26), .Z(
        mux_b[8]) );
  LVT_AO22HSV0 U37 ( .A1(mux_bq[7]), .A2(n35), .B1(b_out[7]), .B2(n26), .Z(
        mux_b[7]) );
  LVT_AO22HSV0 U38 ( .A1(mux_bq[6]), .A2(n35), .B1(b_out[6]), .B2(n26), .Z(
        mux_b[6]) );
  LVT_AO22HSV0 U39 ( .A1(mux_bq[5]), .A2(n35), .B1(b_out[5]), .B2(n26), .Z(
        mux_b[5]) );
  LVT_AO22HSV0 U40 ( .A1(mux_bq[4]), .A2(n35), .B1(b_out[4]), .B2(n26), .Z(
        mux_b[4]) );
  LVT_AO22HSV0 U41 ( .A1(mux_bq[3]), .A2(n35), .B1(b_out[3]), .B2(n26), .Z(
        mux_b[3]) );
  LVT_AO22HSV0 U42 ( .A1(mux_bq[31]), .A2(n35), .B1(b_out[31]), .B2(n26), .Z(
        mux_b[31]) );
  LVT_AO22HSV0 U43 ( .A1(mux_bq[30]), .A2(n35), .B1(b_out[30]), .B2(n26), .Z(
        mux_b[30]) );
  LVT_AO22HSV0 U44 ( .A1(mux_bq[2]), .A2(n35), .B1(b_out[2]), .B2(n26), .Z(
        mux_b[2]) );
  LVT_AO22HSV0 U45 ( .A1(mux_bq[29]), .A2(n35), .B1(b_out[29]), .B2(n26), .Z(
        mux_b[29]) );
  LVT_AO22HSV0 U46 ( .A1(mux_bq[28]), .A2(n35), .B1(b_out[28]), .B2(n26), .Z(
        mux_b[28]) );
  LVT_AO22HSV0 U47 ( .A1(mux_bq[27]), .A2(n35), .B1(b_out[27]), .B2(n26), .Z(
        mux_b[27]) );
  LVT_AO22HSV0 U48 ( .A1(mux_bq[26]), .A2(n35), .B1(b_out[26]), .B2(n26), .Z(
        mux_b[26]) );
  LVT_AO22HSV0 U49 ( .A1(mux_bq[25]), .A2(n35), .B1(b_out[25]), .B2(n26), .Z(
        mux_b[25]) );
  LVT_AO22HSV0 U50 ( .A1(mux_bq[24]), .A2(n35), .B1(b_out[24]), .B2(n26), .Z(
        mux_b[24]) );
  LVT_AO22HSV0 U51 ( .A1(mux_bq[23]), .A2(n35), .B1(b_out[23]), .B2(n26), .Z(
        mux_b[23]) );
  LVT_AO22HSV0 U52 ( .A1(mux_bq[22]), .A2(n35), .B1(b_out[22]), .B2(n26), .Z(
        mux_b[22]) );
  LVT_AO22HSV0 U53 ( .A1(mux_bq[21]), .A2(n35), .B1(b_out[21]), .B2(n26), .Z(
        mux_b[21]) );
  LVT_AO22HSV0 U54 ( .A1(mux_bq[20]), .A2(n35), .B1(b_out[20]), .B2(n26), .Z(
        mux_b[20]) );
  LVT_AO22HSV0 U55 ( .A1(mux_bq[1]), .A2(n35), .B1(b_out[1]), .B2(n26), .Z(
        mux_b[1]) );
  LVT_AO22HSV0 U56 ( .A1(mux_bq[19]), .A2(n35), .B1(b_out[19]), .B2(n26), .Z(
        mux_b[19]) );
  LVT_AO22HSV0 U57 ( .A1(mux_bq[18]), .A2(n35), .B1(b_out[18]), .B2(n26), .Z(
        mux_b[18]) );
  LVT_AO22HSV0 U58 ( .A1(mux_bq[17]), .A2(n35), .B1(b_out[17]), .B2(n26), .Z(
        mux_b[17]) );
  LVT_AO22HSV0 U59 ( .A1(mux_bq[16]), .A2(n35), .B1(b_out[16]), .B2(n26), .Z(
        mux_b[16]) );
  LVT_AO22HSV0 U60 ( .A1(mux_bq[15]), .A2(n35), .B1(b_out[15]), .B2(n26), .Z(
        mux_b[15]) );
  LVT_AO22HSV0 U61 ( .A1(mux_bq[14]), .A2(n35), .B1(b_out[14]), .B2(n26), .Z(
        mux_b[14]) );
  LVT_AO22HSV0 U62 ( .A1(mux_bq[13]), .A2(n35), .B1(b_out[13]), .B2(n26), .Z(
        mux_b[13]) );
  LVT_AO22HSV0 U63 ( .A1(mux_bq[12]), .A2(n35), .B1(b_out[12]), .B2(n26), .Z(
        mux_b[12]) );
  LVT_AO22HSV0 U64 ( .A1(mux_bq[11]), .A2(n35), .B1(b_out[11]), .B2(n26), .Z(
        mux_b[11]) );
  LVT_AO22HSV0 U65 ( .A1(mux_bq[10]), .A2(n35), .B1(b_out[10]), .B2(n26), .Z(
        mux_b[10]) );
  LVT_AO22HSV0 U66 ( .A1(mux_bq[0]), .A2(n35), .B1(b_out[0]), .B2(n26), .Z(
        mux_b[0]) );
  LVT_AOI21HSV0 U69 ( .A1(n4), .A2(n5), .B(n26), .ZN(\c_t_i_1_in[0] ) );
  LVT_AND4HSV0 U71 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .Z(n5) );
  LVT_NOR4HSV0 U72 ( .A1(l_t_i_1_in[9]), .A2(l_t_i_1_in[8]), .A3(l_t_i_1_in[7]), .A4(l_t_i_1_in[6]), .ZN(n9) );
  LVT_NOR4HSV0 U73 ( .A1(l_t_i_1_in[5]), .A2(l_t_i_1_in[4]), .A3(l_t_i_1_in[3]), .A4(l_t_i_1_in[30]), .ZN(n8) );
  LVT_NOR4HSV0 U74 ( .A1(l_t_i_1_in[2]), .A2(l_t_i_1_in[29]), .A3(
        l_t_i_1_in[28]), .A4(l_t_i_1_in[27]), .ZN(n7) );
  LVT_NOR4HSV0 U75 ( .A1(l_t_i_1_in[26]), .A2(l_t_i_1_in[25]), .A3(
        l_t_i_1_in[24]), .A4(l_t_i_1_in[23]), .ZN(n6) );
  LVT_AND4HSV0 U76 ( .A1(n10), .A2(n11), .A3(n12), .A4(n13), .Z(n4) );
  LVT_NOR4HSV0 U77 ( .A1(l_t_i_1_in[22]), .A2(l_t_i_1_in[21]), .A3(
        l_t_i_1_in[20]), .A4(l_t_i_1_in[1]), .ZN(n13) );
  LVT_NOR4HSV0 U78 ( .A1(l_t_i_1_in[19]), .A2(l_t_i_1_in[18]), .A3(
        l_t_i_1_in[17]), .A4(l_t_i_1_in[16]), .ZN(n12) );
  LVT_NOR4HSV0 U79 ( .A1(l_t_i_1_in[15]), .A2(l_t_i_1_in[14]), .A3(
        l_t_i_1_in[13]), .A4(l_t_i_1_in[12]), .ZN(n11) );
  LVT_NOR3HSV0 U80 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[11]), .A3(
        l_t_i_1_in[10]), .ZN(n10) );
  regist_32bit_35 u0 ( .clk(clk), .rstn(n78), .in(a_in), .out(l_a) );
  regist_32bit_34 u1 ( .clk(clk), .rstn(n78), .in(b_in), .out(b_out) );
  regist_32bit_33 u2 ( .clk(clk), .rstn(n78), .in(g_in), .out(l_g) );
  regist_1bit_23 u3 ( .clk(clk), .rstn(n78), .in(ctr), .out(l_ctr) );
  regist_1bit_22 u4 ( .clk(clk), .rstn(n78), .in(n35), .out(ctro) );
  regist_31bit_23 u5 ( .clk(clk), .rstn(n78), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_31bit_22 u6 ( .clk(clk), .rstn(n78), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_21 u7 ( .clk(clk), .rstn(n78), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_32bit_32 u9 ( .clk(clk), .rstn(n78), .in(mux_b), .out(mux_bq) );
  regist_1bit_20 u10 ( .clk(clk), .rstn(n78), .in(to_1), .out(ti_1) );
  regist_31bit_21 u11 ( .clk(clk), .rstn(n78), .in({n75, n65, to_7[28:21], n57, 
        to_7[19], n58, n59, to_7[16:15], n71, n72, to_7[12], n24, to_7[10], 
        n60, to_7[8:6], n61, n62, to_7[3], n63, n73, n74}), .out(ti_7) );
  PE_core_5 pe ( .a_in(l_a), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, n75, 
        n65, to_7[28:21], n57, to_7[19], n58, n59, to_7[16:15], n71, n72, 
        to_7[12], n24, to_7[10], n60, to_7[8:6], n61, n62, to_7[3], n63, n73, 
        n74}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(go), 
        .t_i_1_out(to), .t_i_2_out({t_i_2_out[30:27], n80, t_i_2_out[25:0]}), 
        .t_i_1_out_0(t_i_1_out_0) );
  regist_32bit_31 u12 ( .clk(clk), .rstn(n78), .in(ao), .out(a_out) );
  regist_32bit_30 u13 ( .clk(clk), .rstn(n78), .in(go), .out(g_out) );
  regist_31bit_20 u14 ( .clk(clk), .rstn(n78), .in(to), .out(t_i_1_out) );
  LVT_INHSV8 U2 ( .I(n43), .ZN(n73) );
  LVT_NAND2HSV4 U3 ( .A1(n14), .A2(n15), .ZN(to_7[27]) );
  LVT_INHSV5 U4 ( .I(n53), .ZN(n60) );
  LVT_INHSV10 U5 ( .I(n40), .ZN(n74) );
  LVT_INHSV4 U6 ( .I(n48), .ZN(n72) );
  LVT_AOI22HSV2 U7 ( .A1(ti_7[4]), .A2(ctro), .B1(t_i_2_out[4]), .B2(n1), .ZN(
        n52) );
  LVT_INHSV4 U8 ( .I(n27), .ZN(n63) );
  LVT_NAND2HSV4 U9 ( .A1(n47), .A2(n46), .ZN(to_7[7]) );
  LVT_NAND2HSV4 U10 ( .A1(n68), .A2(n69), .ZN(to_7[12]) );
  LVT_IAO22HSV4 U11 ( .B1(t_i_2_out[2]), .B2(n1), .A1(n28), .A2(n1), .ZN(n27)
         );
  LVT_CLKNHSV6 U12 ( .I(l_ctr), .ZN(n3) );
  LVT_INHSV4 U13 ( .I(n64), .ZN(n75) );
  LVT_CLKNAND2HSV8 U14 ( .A1(l_t_i_1_in_0), .A2(n3), .ZN(n77) );
  LVT_AOI22HSV4 U15 ( .A1(ti_7[13]), .A2(ctro), .B1(t_i_2_out[13]), .B2(n1), 
        .ZN(n48) );
  LVT_NAND2HSV8 U16 ( .A1(n39), .A2(n38), .ZN(to_7[25]) );
  LVT_NAND2HSV4 U17 ( .A1(ti_1), .A2(l_ctr), .ZN(n76) );
  LVT_NAND2HSV8 U18 ( .A1(n37), .A2(n36), .ZN(to_7[8]) );
  LVT_NAND2HSV12 U19 ( .A1(n76), .A2(n77), .ZN(to_1) );
  LVT_CLKNAND2HSV8 U20 ( .A1(n22), .A2(n23), .ZN(to_7[3]) );
  LVT_IAO22HSV4 U21 ( .B1(t_i_2_out[14]), .B2(n1), .A1(n31), .A2(n1), .ZN(n30)
         );
  LVT_NAND2HSV4 U22 ( .A1(n44), .A2(n45), .ZN(to_7[24]) );
  LVT_NAND2HSV4 U23 ( .A1(t_i_2_out[25]), .A2(n1), .ZN(n39) );
  LVT_NAND2HSV4 U24 ( .A1(t_i_2_out[12]), .A2(n1), .ZN(n69) );
  LVT_NAND2HSV8 U25 ( .A1(n41), .A2(n42), .ZN(to_7[21]) );
  LVT_INHSV4SR U26 ( .I(n54), .ZN(n61) );
  LVT_INHSV6SR U27 ( .I(n50), .ZN(n57) );
  LVT_INHSV4 U28 ( .I(n30), .ZN(n71) );
  LVT_CLKNAND2HSV3 U29 ( .A1(n16), .A2(n17), .ZN(to_7[19]) );
  LVT_INHSV4SR U30 ( .I(n52), .ZN(n62) );
  LVT_CLKNAND2HSV4 U31 ( .A1(n25), .A2(n29), .ZN(to_7[22]) );
  LVT_CLKNAND2HSV3 U32 ( .A1(t_i_2_out[22]), .A2(n1), .ZN(n29) );
  LVT_IAO22HSV0 U33 ( .B1(t_i_2_out[18]), .B2(n1), .A1(n33), .A2(n1), .ZN(n32)
         );
  LVT_NAND2HSV0P5 U34 ( .A1(ti_7[27]), .A2(ctro), .ZN(n14) );
  LVT_CLKNAND2HSV3 U67 ( .A1(t_i_2_out[27]), .A2(n1), .ZN(n15) );
  LVT_NAND2HSV0 U68 ( .A1(ti_7[19]), .A2(ctro), .ZN(n16) );
  LVT_CLKNAND2HSV4 U70 ( .A1(t_i_2_out[19]), .A2(n1), .ZN(n17) );
  LVT_INHSV10 U81 ( .I(n49), .ZN(n65) );
  LVT_CLKNAND2HSV8 U82 ( .A1(n20), .A2(n21), .ZN(to_7[10]) );
  LVT_NAND2HSV4 U83 ( .A1(t_i_2_out[10]), .A2(n1), .ZN(n21) );
  LVT_INHSV2 U84 ( .I(n32), .ZN(n58) );
  LVT_CLKNAND2HSV2 U85 ( .A1(t_i_2_out[24]), .A2(n1), .ZN(n45) );
  LVT_NAND2HSV4 U86 ( .A1(t_i_2_out[28]), .A2(n1), .ZN(n56) );
  LVT_INHSV6 U87 ( .I(ctro), .ZN(n1) );
  LVT_INHSV2 U88 ( .I(ti_7[2]), .ZN(n28) );
  LVT_CLKNHSV4 U89 ( .I(n79), .ZN(n78) );
  LVT_NAND2HSV2 U90 ( .A1(ti_7[23]), .A2(ctro), .ZN(n18) );
  LVT_CLKNAND2HSV3 U91 ( .A1(t_i_2_out[23]), .A2(n1), .ZN(n19) );
  LVT_CLKNAND2HSV8 U92 ( .A1(n18), .A2(n19), .ZN(to_7[23]) );
  LVT_NAND2HSV2 U93 ( .A1(ti_7[10]), .A2(ctro), .ZN(n20) );
  LVT_NAND2HSV2 U94 ( .A1(ti_7[3]), .A2(ctro), .ZN(n22) );
  LVT_CLKNAND2HSV3 U95 ( .A1(t_i_2_out[3]), .A2(n1), .ZN(n23) );
  LVT_NAND2HSV4 U96 ( .A1(t_i_2_out[7]), .A2(n1), .ZN(n47) );
  LVT_AO22HSV4 U97 ( .A1(ti_7[11]), .A2(ctro), .B1(t_i_2_out[11]), .B2(n1), 
        .Z(n24) );
  LVT_INHSV2 U98 ( .I(l_t_i_1_in_0), .ZN(n2) );
  LVT_NAND2HSV2 U99 ( .A1(ti_7[22]), .A2(ctro), .ZN(n25) );
  LVT_INHSV2 U100 ( .I(ti_7[18]), .ZN(n33) );
  LVT_INHSV2 U101 ( .I(ti_7[14]), .ZN(n31) );
  LVT_INHSV2 U102 ( .I(n34), .ZN(n26) );
  LVT_CLKNAND2HSV4 U103 ( .A1(t_i_2_out[8]), .A2(n1), .ZN(n37) );
  LVT_NAND2HSV8 U104 ( .A1(n67), .A2(n66), .ZN(to_7[6]) );
  LVT_CLKNAND2HSV8 U105 ( .A1(t_i_2_out[6]), .A2(n1), .ZN(n67) );
  LVT_CLKNAND2HSV4 U106 ( .A1(t_i_2_out[21]), .A2(n1), .ZN(n42) );
  LVT_INHSV4 U107 ( .I(n51), .ZN(n59) );
  LVT_INHSV0SR U108 ( .I(n3), .ZN(n34) );
  LVT_NOR2HSV0P5 U109 ( .A1(n2), .A2(n26), .ZN(c_t_i_1_in_0) );
  LVT_BUFHSV2RT U110 ( .I(n34), .Z(n35) );
  LVT_NAND2HSV0 U111 ( .A1(ti_7[8]), .A2(ctro), .ZN(n36) );
  LVT_NAND2HSV0 U112 ( .A1(ti_7[25]), .A2(ctro), .ZN(n38) );
  LVT_AO22HSV4 U113 ( .A1(ti_7[16]), .A2(ctro), .B1(t_i_2_out[16]), .B2(n1), 
        .Z(to_7[16]) );
  LVT_AOI22HSV4 U114 ( .A1(ti_7[0]), .A2(ctro), .B1(t_i_2_out[0]), .B2(n1), 
        .ZN(n40) );
  LVT_NAND2HSV0 U115 ( .A1(ti_7[21]), .A2(ctro), .ZN(n41) );
  LVT_AOI22HSV4 U116 ( .A1(ti_7[1]), .A2(ctro), .B1(t_i_2_out[1]), .B2(n1), 
        .ZN(n43) );
  LVT_NAND2HSV0 U117 ( .A1(ti_7[24]), .A2(ctro), .ZN(n44) );
  LVT_NAND2HSV0 U118 ( .A1(ti_7[7]), .A2(ctro), .ZN(n46) );
  LVT_AOI22HSV4 U119 ( .A1(ti_7[29]), .A2(ctro), .B1(t_i_2_out[29]), .B2(n1), 
        .ZN(n49) );
  LVT_AOI22HSV4 U120 ( .A1(ti_7[20]), .A2(ctro), .B1(t_i_2_out[20]), .B2(n1), 
        .ZN(n50) );
  LVT_AOI22HSV4 U121 ( .A1(ti_7[17]), .A2(ctro), .B1(t_i_2_out[17]), .B2(n1), 
        .ZN(n51) );
  LVT_AOI22HSV4 U122 ( .A1(ti_7[9]), .A2(ctro), .B1(t_i_2_out[9]), .B2(n1), 
        .ZN(n53) );
  LVT_AOI22HSV4 U123 ( .A1(ti_7[5]), .A2(ctro), .B1(t_i_2_out[5]), .B2(n1), 
        .ZN(n54) );
  LVT_NAND2HSV0 U124 ( .A1(ti_7[28]), .A2(ctro), .ZN(n55) );
  LVT_CLKNAND2HSV8 U125 ( .A1(n55), .A2(n56), .ZN(to_7[28]) );
  LVT_AOI22HSV4 U126 ( .A1(ti_7[30]), .A2(ctro), .B1(t_i_2_out[30]), .B2(n1), 
        .ZN(n64) );
  LVT_NAND2HSV0 U127 ( .A1(ti_7[6]), .A2(ctro), .ZN(n66) );
  LVT_NAND2HSV0 U128 ( .A1(ti_7[12]), .A2(ctro), .ZN(n68) );
  LVT_BUFHSV2RT U129 ( .I(n80), .Z(t_i_2_out[26]) );
  LVT_AO22HSV4 U130 ( .A1(ti_7[15]), .A2(ctro), .B1(t_i_2_out[15]), .B2(n1), 
        .Z(to_7[15]) );
  LVT_AO22HSV4 U131 ( .A1(ti_7[26]), .A2(ctro), .B1(n80), .B2(n1), .Z(to_7[26]) );
  LVT_INHSV2 U132 ( .I(rstn), .ZN(n79) );
endmodule


module regist_32bit_29 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3, n4;

  LVT_DRNQHSV4 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV4 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV4 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV4 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n3), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n3), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n3), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n3), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n3), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n3), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n3), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n3), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_INHSV2 U3 ( .I(n4), .ZN(n2) );
  LVT_INHSV2 U4 ( .I(n4), .ZN(n1) );
  LVT_INHSV2 U5 ( .I(rstn), .ZN(n4) );
  LVT_INHSV2 U6 ( .I(n4), .ZN(n3) );
endmodule


module regist_32bit_28 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3, n4;

  LVT_DRNQHSV2 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n3), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n3), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n3), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n3), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n3), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n3), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n3), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n3), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n4) );
  LVT_INHSV2 U4 ( .I(n4), .ZN(n3) );
  LVT_INHSV2 U5 ( .I(n4), .ZN(n2) );
  LVT_INHSV2 U6 ( .I(n4), .ZN(n1) );
endmodule


module regist_32bit_27 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n7, n1, n3, n4, n5, n6;

  LVT_DRNQHSV4 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n3), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n5), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n3), .Q(out[31]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n3), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n3), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n3), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n3), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n4), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n4), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n4), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n4), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n4), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n4), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n4), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n4), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n4), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n4), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n4), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n4), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n5), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n5), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n5), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n5), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n5), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n5), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n5), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n3), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n3), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n3), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n3), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n3), .Q(n7) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n3), .Q(out[29]) );
  LVT_CLKNHSV4 U3 ( .I(n1), .ZN(out[27]) );
  LVT_INHSV2 U4 ( .I(n7), .ZN(n1) );
  LVT_INHSV2 U5 ( .I(n6), .ZN(n4) );
  LVT_INHSV2 U6 ( .I(n6), .ZN(n3) );
  LVT_INHSV2 U7 ( .I(rstn), .ZN(n6) );
  LVT_INHSV2 U8 ( .I(n6), .ZN(n5) );
endmodule


module regist_1bit_19 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;
  wire   n3, n1;

  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(n3) );
  LVT_INHSV20 U3 ( .I(n1), .ZN(out) );
  LVT_INHSV8 U4 ( .I(n3), .ZN(n1) );
endmodule


module regist_1bit_18 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_31bit_19 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2, n3, n4;

  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n1), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n2), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n3), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n3), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n3), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n3), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n3), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n3), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n3), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(n4), .ZN(n2) );
  LVT_INHSV2 U4 ( .I(n4), .ZN(n1) );
  LVT_INHSV2 U5 ( .I(rstn), .ZN(n4) );
  LVT_INHSV2 U6 ( .I(n4), .ZN(n3) );
endmodule


module regist_31bit_18 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n2), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n2), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n1), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n2), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n2), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(rstn), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(rstn), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n1), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n1), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n2), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n2), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n1), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(rstn), .Q(out[11])
         );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n1), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n1), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n2), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n2), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n2), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n2), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n1), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n2), .Q(out[7]) );
  LVT_INHSV2 U3 ( .I(n3), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n2) );
endmodule


module regist_1bit_17 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_32bit_26 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3, n4;

  LVT_DRNQHSV4 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n3), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n3), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n3), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n2), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n2), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n2), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n2), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n2), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n2), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n3), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n3), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n3), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n3), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n3), .Q(out[12]) );
  LVT_INHSV2 U3 ( .I(n4), .ZN(n2) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n4) );
  LVT_INHSV2 U5 ( .I(n4), .ZN(n3) );
  LVT_INHSV2 U6 ( .I(n4), .ZN(n1) );
endmodule


module regist_1bit_16 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV1 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_31bit_17 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n2), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n2), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n2), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n2), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n2), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n1) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n2) );
endmodule


module cell_3_4809 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_154 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_153 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_152 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_151 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_150 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_149 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_148 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_147 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_146 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_145 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_144 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_143 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_142 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_141 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_140 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_139 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_138 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_137 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_136 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_135 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKNAND2HSV2 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_134 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_CLKNAND2HSV1 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_133 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_132 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_131 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_4_130 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U3 ( .A1(n5), .A2(n6), .Z(n7) );
endmodule


module cell_4_129 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_128 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U3 ( .A1(n7), .A2(n8), .Z(t_i_out) );
endmodule


module cell_4_127 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_126 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_125 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n2, n5, n6;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n1), .A2(n2), .Z(t_i_out) );
  LVT_XNOR2HSV4 U3 ( .A1(n5), .A2(n6), .ZN(n1) );
  LVT_XNOR2HSV1 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_4_124 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  LVT_INHSV4SR U1 ( .I(n15), .ZN(n8) );
  LVT_CLKNAND2HSV1 U2 ( .A1(n15), .A2(n12), .ZN(n10) );
  LVT_CLKNAND2HSV3 U3 ( .A1(n6), .A2(n7), .ZN(n15) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n1), .A2(n14), .ZN(n7) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n13), .A2(n5), .ZN(n6) );
  LVT_XNOR2HSV1 U6 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n12) );
  LVT_CLKNAND2HSV8 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n13) );
  LVT_CLKNAND2HSV4 U8 ( .A1(n10), .A2(n11), .ZN(t_i_out) );
  LVT_NAND2HSV4 U9 ( .A1(n8), .A2(n9), .ZN(n11) );
  LVT_INHSV4 U10 ( .I(n13), .ZN(n1) );
  LVT_CLKNHSV1 U11 ( .I(n14), .ZN(n5) );
  LVT_NAND2HSV0P5 U12 ( .A1(b_in), .A2(a_in), .ZN(n14) );
  LVT_CLKNHSV0P5 U13 ( .I(n12), .ZN(n9) );
endmodule


module row_1_4 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [31:0] t_i_1_in;
  input [30:0] t_i_2_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_3_4809 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_154 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(t_i_1_out[1])
         );
  cell_4_153 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(t_i_1_out[2])
         );
  cell_4_152 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(t_i_1_out[3])
         );
  cell_4_151 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(t_i_1_out[4])
         );
  cell_4_150 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(t_i_1_out[5])
         );
  cell_4_149 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(t_i_1_out[6])
         );
  cell_4_148 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(t_i_1_out[7])
         );
  cell_4_147 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_2_in(t_i_2_in[7]), .t_i_out(t_i_1_out[8])
         );
  cell_4_146 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[9]), .t_i_2_in(t_i_2_in[8]), .t_i_out(t_i_1_out[9])
         );
  cell_4_145 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[10]), .t_i_2_in(t_i_2_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_4_144 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[11]), .t_i_2_in(t_i_2_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_4_143 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[12]), .t_i_2_in(t_i_2_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_4_142 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[13]), .t_i_2_in(t_i_2_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_4_141 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[14]), .t_i_2_in(t_i_2_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_4_140 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[15]), .t_i_2_in(t_i_2_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_4_139 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[16]), .t_i_2_in(t_i_2_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_4_138 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[17]), .t_i_2_in(t_i_2_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_4_137 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[18]), .t_i_2_in(t_i_2_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_4_136 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[19]), .t_i_2_in(t_i_2_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_4_135 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[20]), .t_i_2_in(t_i_2_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_4_134 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[21]), .t_i_2_in(t_i_2_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_4_133 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_2_in(t_i_2_in[21]), .t_i_out(
        t_i_1_out[22]) );
  cell_4_132 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_2_in(t_i_2_in[22]), .t_i_out(
        t_i_1_out[23]) );
  cell_4_131 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_2_in(t_i_2_in[23]), .t_i_out(
        t_i_1_out[24]) );
  cell_4_130 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_2_in(t_i_2_in[24]), .t_i_out(
        t_i_1_out[25]) );
  cell_4_129 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_2_in(t_i_2_in[25]), .t_i_out(
        t_i_1_out[26]) );
  cell_4_128 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_2_in(t_i_2_in[26]), .t_i_out(
        t_i_1_out[27]) );
  cell_4_127 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_2_in(t_i_2_in[27]), .t_i_out(
        t_i_1_out[28]) );
  cell_4_126 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_2_in(t_i_2_in[28]), .t_i_out(
        t_i_1_out[29]) );
  cell_4_125 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_2_in(t_i_2_in[29]), .t_i_out(
        t_i_1_out[30]) );
  cell_4_124 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[31]), .t_i_2_in(t_i_2_in[30]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV2SR U1 ( .I(t_m_1_in), .ZN(n3) );
  LVT_INHSV4 U2 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U3 ( .I(n3), .ZN(n1) );
  LVT_BUFHSV2RT U4 ( .I(n2), .Z(n4) );
endmodule


module cell_2_154 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4808 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4807 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4806 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4805 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4804 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4803 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4802 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4801 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4800 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4799 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4798 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4797 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4796 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4795 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4794 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4793 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4792 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4791 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4790 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4789 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4788 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4787 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4786 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4785 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4784 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4783 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4782 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4781 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4780 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U2 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_4779 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_XNOR2HSV1 U1 ( .A1(t_i_1_in), .A2(n5), .ZN(n4) );
  LVT_OAI21HSV2 U2 ( .A1(n6), .A2(n4), .B(n2), .ZN(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U5 ( .A1(n6), .A2(n4), .ZN(n2) );
endmodule


module cell_3_4778 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV1 U1 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2 U2 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U4 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNAND2HSV3 U5 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV4SR U6 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV8 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV4 U8 ( .A1(n2), .A2(n4), .ZN(n6) );
endmodule


module row_other_154 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_154 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4808 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4807 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4806 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4805 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4804 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4803 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4802 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4801 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4800 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4799 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4798 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4797 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4796 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4795 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4794 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4793 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4792 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4791 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4790 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4789 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4788 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4787 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4786 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4785 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4784 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4783 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4782 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4781 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4780 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4779 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4778 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_153 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4777 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4776 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4775 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4774 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4773 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4772 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4771 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4770 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4769 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4768 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4767 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4766 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4765 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4764 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4763 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV0 U5 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_4762 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4761 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4760 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4759 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4758 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4757 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4756 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4755 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4754 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4753 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4752 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4751 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4750 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_XOR2HSV4 U1 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_CLKAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .Z(n3) );
  LVT_XNOR2HSV4 U3 ( .A1(n3), .A2(t_i_1_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_4749 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV4 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4748 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4747 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0 U1 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV3SR U2 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV4 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U6 ( .A1(n4), .A2(n2), .ZN(n6) );
  LVT_INHSV2 U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_153 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_2_153 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4777 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4776 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4775 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4774 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4773 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4772 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4771 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4770 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4769 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4768 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4767 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4766 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4765 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4764 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4763 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4762 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4761 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4760 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4759 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4758 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4757 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4756 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4755 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4754 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4753 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4752 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4751 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4750 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4749 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4748 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4747 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV3SR U1 ( .I(n2), .ZN(n3) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n2) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n4) );
  LVT_INHSV2 U4 ( .I(n2), .ZN(n1) );
endmodule


module cell_2_152 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4746 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4745 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4744 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4743 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4742 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4741 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4740 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4739 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4738 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4737 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4736 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4735 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4734 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4733 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4732 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4731 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4730 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4729 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4728 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4727 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4726 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4725 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4724 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4723 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4722 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4721 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4720 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4719 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n5), .A2(n6), .Z(t_i_out) );
endmodule


module cell_3_4718 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_4717 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4716 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV4 U1 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV4SR U2 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV1 U4 ( .A1(n7), .A2(n9), .ZN(n5) );
  LVT_NAND2HSV4 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV2SR U6 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV2 U7 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_152 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_152 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4746 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4745 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4744 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4743 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4742 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4741 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4740 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4739 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4738 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4737 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4736 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4735 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4734 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4733 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4732 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4731 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4730 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4729 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4728 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4727 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4726 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4725 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4724 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4723 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4722 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4721 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4720 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4719 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4718 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4717 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4716 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV4 U1 ( .I(n2), .ZN(n1) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n2) );
endmodule


module cell_2_151 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4715 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4714 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4713 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4712 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4711 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4710 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4709 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4708 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4707 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4706 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4705 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4704 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4703 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4702 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4701 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4700 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4699 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4698 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4697 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4696 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4695 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4694 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4693 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4692 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4691 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4690 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4689 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4688 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U2 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_4687 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4686 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_4685 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5, n6, n7, n8, n9;

  LVT_INHSV2SR U1 ( .I(n8), .ZN(n4) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n3), .A2(n8), .ZN(n6) );
  LVT_CLKNAND2HSV1 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV0P5 U4 ( .A1(n9), .A2(n4), .ZN(n5) );
  LVT_CLKNAND2HSV3 U5 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV2 U6 ( .I(n9), .ZN(n3) );
  LVT_CLKAND2HSV2 U7 ( .A1(b_in), .A2(a_in), .Z(n7) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n7), .ZN(n8) );
endmodule


module row_other_151 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_151 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4715 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4714 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4713 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4712 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4711 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4710 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4709 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4708 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4707 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4706 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4705 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4704 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4703 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4702 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4701 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4700 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4699 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4698 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4697 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4696 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4695 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4694 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4693 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4692 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4691 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4690 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4689 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4688 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4687 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4686 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4685 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV4 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_150 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4684 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4683 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4682 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4681 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4680 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4679 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4678 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4677 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4676 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4675 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4674 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4673 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4672 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4671 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4670 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4669 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4668 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4667 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4666 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4665 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4664 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4663 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4662 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4661 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4660 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4659 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_4658 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4657 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4656 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_4655 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4654 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_150 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4, n5;

  cell_2_150 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4684 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4683 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4682 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4681 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4680 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4679 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4678 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4677 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4676 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4675 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4674 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4673 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4672 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4671 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4670 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4669 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4668 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4667 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4666 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4665 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4664 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4663 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4662 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4661 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4660 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4659 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4658 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4657 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4656 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4655 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4654 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV4 U1 ( .I(n3), .ZN(n4) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n3) );
  LVT_INHSV0SR U3 ( .I(t_m_1_in), .ZN(n1) );
  LVT_CLKNHSV0P5 U4 ( .I(n1), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n1), .ZN(n5) );
endmodule


module cell_2_149 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4653 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4652 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4651 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4650 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4649 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4648 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4647 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4646 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4645 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4644 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4643 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4642 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4641 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4640 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4639 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4638 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4637 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4636 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4635 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4634 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4633 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4632 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4631 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4630 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4629 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4628 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4627 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_4626 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4625 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_XOR2HSV0 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U5 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_3_4624 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4623 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U4 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2SR U6 ( .I(n7), .ZN(n4) );
  LVT_INHSV2SR U7 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV2 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
endmodule


module row_other_149 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_149 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4653 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4652 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4651 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4650 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4649 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4648 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4647 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4646 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4645 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4644 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4643 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4642 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4641 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4640 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4639 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4638 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4637 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4636 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4635 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4634 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4633 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4632 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4631 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4630 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4629 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4628 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4627 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4626 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4625 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4624 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4623 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV4 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_148 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4622 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4621 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4620 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4619 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4618 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4617 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4616 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4615 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4614 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4613 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4612 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4611 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4610 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4609 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4608 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4607 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4606 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4605 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4604 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4603 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4602 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4601 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4600 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4599 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4598 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4597 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4596 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4595 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4594 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4593 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4592 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;

  LVT_CLKNHSV2P5 U1 ( .I(n11), .ZN(n2) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n11) );
  LVT_NAND2HSV2 U3 ( .A1(n8), .A2(n9), .ZN(n10) );
  LVT_CLKNHSV2 U4 ( .I(n10), .ZN(n3) );
  LVT_CLKNHSV1 U5 ( .I(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV0P5 U6 ( .A1(n11), .A2(n10), .ZN(n4) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n2), .A2(n3), .ZN(n5) );
  LVT_CLKNAND2HSV3 U8 ( .A1(n4), .A2(n5), .ZN(t_i_out) );
  LVT_CLKAND2HSV2 U9 ( .A1(b_in), .A2(a_in), .Z(n6) );
  LVT_INAND2HSV0 U10 ( .A1(n6), .B1(t_i_1_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U11 ( .A1(n6), .A2(n7), .ZN(n9) );
endmodule


module row_other_148 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_148 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4622 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4621 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4620 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4619 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4618 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4617 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4616 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4615 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4614 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4613 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4612 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4611 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4610 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4609 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4608 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4607 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4606 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4605 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4604 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4603 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4602 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4601 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4600 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4599 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4598 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4597 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4596 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4595 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4594 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4593 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4592 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV4 U1 ( .I(n1), .ZN(n2) );
  LVT_CLKNHSV0 U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_147 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_4591 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4590 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4589 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4588 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4587 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4586 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4585 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4584 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4583 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4582 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4581 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4580 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4579 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4578 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4577 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4576 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4575 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4574 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4573 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4572 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4571 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4570 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4569 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4568 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4567 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4566 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4565 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4564 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4563 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_4562 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module cell_3_4561 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKNAND2HSV1 U2 ( .A1(n6), .A2(n4), .ZN(n2) );
  LVT_OAI21HSV2 U4 ( .A1(n6), .A2(n4), .B(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U5 ( .A1(n5), .A2(t_i_1_in), .ZN(n4) );
endmodule


module row_other_147 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_147 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_4591 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4590 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4589 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4588 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4587 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4586 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4585 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4584 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4583 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4582 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4581 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4580 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4579 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4578 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4577 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4576 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4575 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4574 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4573 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4572 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4571 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4570 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4569 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4568 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4567 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4566 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4565 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4564 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4563 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4562 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4561 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV2 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_146 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_4560 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4559 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4558 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4557 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4556 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4555 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4554 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4553 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4552 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4551 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4550 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4549 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4548 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4547 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4546 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4545 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4544 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4543 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4542 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4541 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4540 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4539 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4538 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4537 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4536 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4535 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4534 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_4533 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4532 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4531 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4530 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_146 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_146 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4560 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4559 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4558 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4557 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4556 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4555 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4554 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4553 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4552 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4551 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4550 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4549 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4548 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4547 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4546 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4545 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4544 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4543 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4542 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4541 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4540 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4539 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4538 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4537 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4536 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4535 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4534 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4533 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4532 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4531 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4530 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV1 U1 ( .I(t_m_1_in), .ZN(n2) );
  LVT_CLKNHSV6 U2 ( .I(n2), .ZN(n1) );
endmodule


module cell_2_145 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4529 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4528 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4527 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4526 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4525 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4524 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4523 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4522 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4521 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4520 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4519 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4518 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4517 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4516 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4515 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4514 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4513 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4512 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4511 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4510 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4509 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4508 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4507 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4506 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4505 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4504 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4503 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4502 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_XOR2HSV2 U2 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_NAND2HSV0P5 U4 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_NAND2HSV2 U6 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV2SR U7 ( .I(n10), .ZN(n4) );
  LVT_INHSV0SR U8 ( .I(n9), .ZN(n5) );
endmodule


module cell_3_4501 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_XOR2HSV0 U1 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0P5 U3 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_CLKNHSV0 U5 ( .I(n8), .ZN(n4) );
  LVT_CLKNHSV2 U6 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV0 U7 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_4500 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4499 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV4 U1 ( .A1(n2), .A2(n4), .ZN(n5) );
  LVT_CLKNAND2HSV2 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV2P5 U4 ( .I(n9), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U6 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNAND2HSV3 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV0P5 U8 ( .A1(n9), .A2(n7), .ZN(n6) );
endmodule


module row_other_145 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_145 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4529 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4528 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4527 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4526 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4525 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4524 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4523 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4522 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4521 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4520 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4519 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4518 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4517 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4516 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4515 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4514 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4513 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4512 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4511 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4510 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4509 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4508 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4507 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4506 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4505 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4504 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4503 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4502 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4501 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4500 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4499 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV8 U1 ( .I(n2), .ZN(n3) );
  LVT_INHSV4SR U2 ( .I(t_m_1_in), .ZN(n2) );
  LVT_BUFHSV4RQ U3 ( .I(n3), .Z(n1) );
endmodule


module cell_2_144 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4498 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4497 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4496 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4495 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4494 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4493 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4492 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4491 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4490 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4489 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4488 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4487 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4486 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4485 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4484 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4483 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4482 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4481 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4480 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4479 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4478 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4477 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4476 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4475 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4474 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4473 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4472 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4471 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4470 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4469 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4468 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;

  LVT_CLKNAND2HSV2 U1 ( .A1(n7), .A2(n8), .ZN(n10) );
  LVT_CLKNAND2HSV1 U2 ( .A1(n10), .A2(n9), .ZN(t_i_out) );
  LVT_NAND2HSV2 U3 ( .A1(n12), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV2 U5 ( .A1(n5), .A2(n6), .ZN(n11) );
  LVT_CLKNHSV2P5 U6 ( .I(n12), .ZN(n2) );
  LVT_INHSV4 U7 ( .I(t_i_1_in), .ZN(n4) );
  LVT_NAND2HSV0 U8 ( .A1(b_in), .A2(a_in), .ZN(n12) );
  LVT_NAND2HSV0 U9 ( .A1(n13), .A2(n11), .ZN(n9) );
  LVT_INHSV1SR U10 ( .I(n13), .ZN(n7) );
  LVT_NAND2HSV1 U11 ( .A1(t_m_1_in), .A2(g_in), .ZN(n13) );
  LVT_INHSV2SR U12 ( .I(n11), .ZN(n8) );
endmodule


module row_other_144 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_144 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4498 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4497 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4496 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4495 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4494 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4493 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4492 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4491 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4490 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4489 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4488 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4487 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4486 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4485 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4484 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4483 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4482 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4481 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4480 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4479 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4478 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4477 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4476 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4475 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4474 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4473 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4472 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4471 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4470 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4469 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4468 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV12SR U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV4SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_143 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4467 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4466 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4465 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4464 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4463 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4462 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4461 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4460 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4459 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4458 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4457 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4456 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4455 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4454 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4453 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4452 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4451 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4450 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4449 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4448 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4447 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4446 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4445 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4444 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4443 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4442 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4441 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4440 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_4439 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4438 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4437 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_143 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_143 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4467 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4466 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4465 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4464 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4463 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4462 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4461 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4460 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4459 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4458 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4457 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4456 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4455 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4454 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4453 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4452 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4451 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4450 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4449 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4448 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4447 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4446 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4445 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4444 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4443 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4442 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4441 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4440 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4439 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4438 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4437 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV6 U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_CLKNHSV12 U2 ( .I(n1), .ZN(n3) );
  LVT_INHSV4SR U3 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_142 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4436 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4435 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4434 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4433 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4432 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4431 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4430 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4429 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4428 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4427 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4426 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4425 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4424 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4423 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4422 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4421 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4420 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4419 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4418 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4417 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4416 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4415 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4414 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4413 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4412 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4411 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4410 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4409 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4408 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4407 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_4406 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKXOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module row_other_142 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_142 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4436 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4435 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4434 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4433 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4432 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4431 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4430 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4429 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4428 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4427 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4426 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4425 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4424 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4423 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4422 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4421 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4420 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4419 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4418 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4417 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4416 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4415 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4414 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4413 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4412 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4411 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4410 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4409 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4408 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4407 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4406 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV2 U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_CLKNHSV10 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_141 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4405 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4404 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4403 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4402 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4401 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4400 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4399 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4398 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4397 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4396 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4395 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4394 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4393 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4392 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4391 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4390 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4389 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4388 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4387 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4386 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4385 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4384 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4383 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4382 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4381 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4380 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4379 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4378 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4377 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4376 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_4375 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_141 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_141 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4405 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4404 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4403 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4402 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4401 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4400 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4399 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4398 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4397 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4396 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4395 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4394 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4393 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4392 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4391 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4390 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4389 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4388 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4387 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4386 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4385 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4384 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4383 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4382 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4381 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4380 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4379 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4378 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4377 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4376 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4375 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV8SR U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV3SR U2 ( .I(t_m_1_in), .ZN(n1) );
  LVT_CLKNHSV0P5 U3 ( .I(n1), .ZN(n3) );
endmodule


module cell_2_140 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_4374 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4373 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4372 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4371 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4370 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4369 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4368 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4367 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4366 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4365 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4364 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4363 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4362 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4361 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4360 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4359 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4358 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4357 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4356 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4355 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4354 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4353 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4352 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4351 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV3 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4350 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4349 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4348 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4347 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4346 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_4345 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV1 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0P5 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U3 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0P5 U4 ( .I(n8), .ZN(n4) );
  LVT_CLKNHSV2 U5 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV8 U6 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV4 U7 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV0 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_4344 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4;

  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n4) );
  LVT_CLKAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .Z(n2) );
  LVT_XNOR2HSV4 U3 ( .A1(n4), .A2(n3), .ZN(t_i_out) );
  LVT_XOR2HSV4 U4 ( .A1(n2), .A2(t_i_1_in), .Z(n3) );
endmodule


module row_other_140 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4, n5;

  cell_2_140 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4374 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4373 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4372 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4371 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4370 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4369 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4368 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4367 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4366 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4365 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4364 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4363 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4362 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4361 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4360 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4359 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4358 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4357 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4356 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4355 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4354 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4353 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4352 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4351 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4350 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4349 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4348 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4347 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4346 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4345 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4344 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV3SR U1 ( .I(n2), .ZN(n3) );
  LVT_INHSV6 U2 ( .I(n4), .ZN(n1) );
  LVT_INHSV0SR U3 ( .I(t_m_1_in), .ZN(n2) );
  LVT_BUFHSV2RT U4 ( .I(n1), .Z(n5) );
  LVT_INHSV0SR U5 ( .I(t_m_1_in), .ZN(n4) );
endmodule


module cell_2_139 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4343 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4342 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4341 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4340 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4339 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4338 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4337 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4336 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4335 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4334 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4333 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4332 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4331 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4330 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4329 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4328 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4327 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4326 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4325 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4324 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4323 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4322 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4321 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4320 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4319 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4318 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4317 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4316 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4315 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4314 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKXOR2HSV2 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U3 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U4 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U5 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_4313 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9, n10;

  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV0P5 U2 ( .A1(n5), .A2(n6), .ZN(n8) );
  LVT_OAI21HSV2 U3 ( .A1(n10), .A2(n8), .B(n7), .ZN(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(n10), .A2(n8), .ZN(n7) );
  LVT_NAND2HSV2 U5 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV0P5 U6 ( .A1(n9), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U7 ( .I(n9), .ZN(n2) );
  LVT_INHSV2 U8 ( .I(t_i_1_in), .ZN(n4) );
  LVT_NAND2HSV0 U9 ( .A1(b_in), .A2(a_in), .ZN(n9) );
endmodule


module row_other_139 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4, n5, n6;

  cell_2_139 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4343 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4342 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4341 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4340 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4339 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4338 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4337 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4336 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4335 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4334 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4333 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4332 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4331 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4330 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4329 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4328 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4327 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4326 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4325 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4324 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n6), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4323 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4322 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n6), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4321 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n6), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4320 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n6), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4319 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n6), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4318 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n6), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4317 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n6), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4316 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n6), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4315 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4314 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4313 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV4 U1 ( .I(t_m_1_in), .ZN(n5) );
  LVT_INHSV0SR U2 ( .I(n6), .ZN(n1) );
  LVT_INHSV2 U3 ( .I(n1), .ZN(n2) );
  LVT_INHSV4SR U4 ( .I(n5), .ZN(n6) );
  LVT_BUFHSV2RT U5 ( .I(n6), .Z(n3) );
  LVT_INHSV0SR U6 ( .I(n5), .ZN(n4) );
endmodule


module cell_2_138 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_4312 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4311 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4310 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4309 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4308 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4307 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4306 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4305 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4304 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4303 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4302 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4301 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4300 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4299 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4298 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4297 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4296 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4295 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4294 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4293 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4292 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4291 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4290 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4289 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4288 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4287 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4286 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4285 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4284 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4283 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4282 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_138 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_138 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4312 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4311 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4310 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4309 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4308 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4307 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4306 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4305 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4304 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4303 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4302 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4301 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4300 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4299 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4298 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4297 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4296 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4295 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4294 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4293 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4292 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4291 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4290 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4289 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4288 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4287 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4286 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4285 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4284 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4283 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4282 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV6RT U1 ( .I(t_m_1_in), .Z(n3) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U3 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_137 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4281 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4280 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4279 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4278 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4277 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4276 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4275 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4274 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4273 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4272 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4271 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4270 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4269 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4268 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4267 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4266 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4265 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4264 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4263 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4262 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4261 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4260 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4259 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4258 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4257 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4256 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4255 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4254 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4253 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV3 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4252 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4251 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_137 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_137 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_4281 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4280 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4279 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4278 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4277 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4276 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4275 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4274 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4273 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4272 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4271 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4270 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4269 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4268 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4267 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4266 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4265 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4264 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4263 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4262 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4261 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4260 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4259 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4258 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4257 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4256 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4255 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4254 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4253 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4252 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4251 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_136 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4250 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4249 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4248 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4247 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4246 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4245 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4244 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4243 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4242 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4241 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4240 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4239 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4238 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4237 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4236 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4235 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4234 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4233 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4232 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4231 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4230 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4229 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4228 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4227 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4226 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4225 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4224 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4223 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4222 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4221 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_4220 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNHSV2P5 U2 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U4 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U8 ( .I(n9), .ZN(n2) );
endmodule


module row_other_136 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_136 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4250 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4249 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4248 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4247 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4246 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4245 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4244 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4243 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4242 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4241 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4240 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4239 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4238 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4237 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4236 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4235 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4234 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4233 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4232 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4231 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4230 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4229 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4228 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4227 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4226 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4225 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4224 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4223 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4222 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4221 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4220 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV8 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV2P5 U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_135 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_4219 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4218 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4217 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4216 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4215 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4214 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4213 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4212 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4211 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4210 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4209 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4208 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4207 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4206 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4205 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4204 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4203 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4202 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4201 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4200 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4199 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4198 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4197 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4196 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4195 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4194 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4193 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4192 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV3 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0P5 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNAND2HSV3 U3 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_CLKNHSV0P5 U4 ( .I(n8), .ZN(n4) );
  LVT_CLKNHSV2P5 U5 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV8 U6 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV2 U7 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV0 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_4191 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4190 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4189 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_CLKNHSV2 U1 ( .I(n6), .ZN(n4) );
  LVT_INHSV2P5 U2 ( .I(n8), .ZN(n2) );
  LVT_NAND2HSV4 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_IOA21HSV2 U5 ( .A1(n8), .A2(n6), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV2 U6 ( .A1(n2), .A2(n4), .ZN(n5) );
  LVT_XNOR2HSV4 U7 ( .A1(n7), .A2(t_i_1_in), .ZN(n6) );
endmodule


module row_other_135 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_135 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4219 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4218 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4217 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4216 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4215 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4214 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4213 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4212 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4211 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4210 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4209 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4208 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4207 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4206 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4205 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4204 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4203 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4202 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4201 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4200 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4199 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4198 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4197 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4196 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4195 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4194 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4193 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4192 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4191 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4190 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4189 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV6 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_134 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_4188 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4187 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4186 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4185 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4184 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4183 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4182 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4181 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4180 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4179 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4178 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4177 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4176 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4175 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4174 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4173 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4172 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4171 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4170 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4169 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4168 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4167 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4166 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4165 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4164 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_NAND2HSV2 U1 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U3 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U5 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_4163 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4162 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_XOR2HSV0 U1 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0 U3 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0SR U5 ( .I(n8), .ZN(n4) );
  LVT_INHSV2 U6 ( .I(t_i_1_in), .ZN(n5) );
  LVT_CLKNAND2HSV4 U7 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_4161 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV2 U1 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_CLKNAND2HSV1 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_CLKNHSV0 U5 ( .I(n10), .ZN(n4) );
  LVT_INHSV4 U6 ( .I(n9), .ZN(n5) );
  LVT_XOR2HSV4 U7 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_NAND2HSV0 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_4160 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4159 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4158 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U1 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV4 U4 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNHSV2P5 U5 ( .I(n9), .ZN(n2) );
  LVT_INHSV2 U6 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV3 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV2 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_134 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_134 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_4188 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4187 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4186 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4185 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4184 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4183 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4182 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4181 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4180 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4179 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4178 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4177 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4176 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4175 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4174 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4173 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4172 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4171 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4170 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4169 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4168 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4167 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4166 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4165 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4164 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4163 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4162 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4161 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4160 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4159 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4158 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV2 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_133 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_4157 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4156 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4155 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4154 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4153 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4152 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4151 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4150 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4149 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4148 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4147 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4146 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4145 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4144 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4143 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4142 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4141 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4140 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4139 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4138 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4137 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4136 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4135 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4134 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4133 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4132 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4131 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4130 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4129 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4128 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4127 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_XNOR2HSV4 U1 ( .A1(n7), .A2(t_i_1_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U2 ( .A1(n8), .A2(n6), .ZN(n4) );
  LVT_INAND2HSV4 U4 ( .A1(n8), .B1(n2), .ZN(n5) );
  LVT_CLKNAND2HSV8 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n5), .A2(n4), .ZN(t_i_out) );
  LVT_INHSV2 U7 ( .I(n6), .ZN(n2) );
endmodule


module row_other_133 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4, n5;

  cell_2_133 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4157 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4156 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4155 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4154 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4153 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4152 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4151 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4150 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4149 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4148 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4147 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4146 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4145 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4144 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4143 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4142 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4141 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4140 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4139 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4138 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4137 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4136 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4135 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4134 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4133 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4132 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4131 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4130 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4129 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4128 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4127 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n4) );
  LVT_CLKNHSV4 U2 ( .I(n3), .ZN(n1) );
  LVT_INHSV2 U3 ( .I(n4), .ZN(n3) );
  LVT_INHSV12SR U4 ( .I(n1), .ZN(n2) );
  LVT_CLKNHSV0P5 U5 ( .I(n4), .ZN(n5) );
endmodule


module cell_2_132 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4126 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4125 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4124 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4123 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4122 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4121 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4120 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4119 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4118 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4117 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4116 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4115 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4114 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4113 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4112 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4111 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4110 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4109 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4108 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4107 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4106 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4105 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4104 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4103 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4102 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4101 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_XOR2HSV0 U1 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV2 U2 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U6 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0SR U7 ( .I(n8), .ZN(n4) );
  LVT_INHSV2 U8 ( .I(t_i_1_in), .ZN(n5) );
endmodule


module cell_3_4100 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4099 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_4098 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4097 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4096 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV3 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV3SR U5 ( .I(n9), .ZN(n2) );
  LVT_INHSV3SR U6 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV4 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_132 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1;

  cell_2_132 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_4126 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4125 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4124 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4123 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4122 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4121 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4120 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4119 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4118 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4117 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4116 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4115 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4114 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4113 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4112 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4111 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4110 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4109 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4108 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4107 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4106 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4105 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4104 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4103 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4102 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4101 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4100 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4099 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4098 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4097 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4096 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV4 U1 ( .I(t_m_1_in), .Z(n1) );
endmodule


module cell_2_131 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_4095 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4094 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4093 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4092 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4091 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4090 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4089 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4088 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4087 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4086 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4085 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4084 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4083 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4082 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4081 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4080 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4079 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4078 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4077 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4076 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4075 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4074 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4073 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4072 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4071 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4070 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4069 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4068 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4067 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4066 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4065 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV2 U1 ( .I(n10), .ZN(n4) );
  LVT_CLKNAND2HSV1 U2 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_INHSV2SR U4 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV2 U5 ( .A1(n7), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U6 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_CLKNAND2HSV3 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_XOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
endmodule


module row_other_131 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_2_131 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4095 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4094 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4093 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4092 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4091 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4090 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4089 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4088 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4087 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4086 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4085 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4084 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4083 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4082 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4081 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4080 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4079 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4078 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4077 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4076 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4075 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4074 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4073 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4072 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4071 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4070 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4069 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4068 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4067 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4066 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4065 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_CLKNHSV6 U2 ( .I(n1), .ZN(n2) );
  LVT_INHSV2SR U3 ( .I(n3), .ZN(n4) );
  LVT_INHSV0SR U4 ( .I(t_m_1_in), .ZN(n3) );
endmodule


module cell_2_130 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4064 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4063 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4062 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4061 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4060 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4059 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4058 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4057 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4056 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4055 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_INHSV0SR U4 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XOR2HSV2 U6 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
endmodule


module cell_3_4054 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4053 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4052 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4051 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4050 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4049 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4048 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4047 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4046 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4045 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4044 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4043 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4042 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4041 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4040 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4039 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4038 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4037 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4036 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4035 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4034 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV2 U1 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(n7), .A2(n9), .ZN(n5) );
  LVT_INHSV0P5SR U4 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_130 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_130 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4064 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4063 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4062 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4061 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4060 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4059 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4058 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4057 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4056 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4055 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4054 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4053 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4052 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4051 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4050 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4049 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4048 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4047 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4046 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4045 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4044 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4043 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4042 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4041 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4040 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4039 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4038 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4037 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4036 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4035 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4034 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV16 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV6 U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_129 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_4033 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4032 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4031 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4030 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4029 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4028 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4027 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4026 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4025 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4024 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4023 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4022 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4021 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4020 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4019 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4018 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4017 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4016 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4015 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4014 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4013 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4012 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4011 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4010 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4009 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4008 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4007 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_4006 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4005 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4004 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4003 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n5), .A2(n9), .ZN(n7) );
  LVT_CLKNAND2HSV3 U3 ( .A1(n7), .A2(n6), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U4 ( .A1(n8), .A2(t_i_1_in), .ZN(n4) );
  LVT_INHSV2 U5 ( .I(n10), .ZN(n5) );
  LVT_NAND2HSV0 U6 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U7 ( .A1(n10), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module row_other_129 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_129 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_4033 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4032 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4031 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_4030 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_4029 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_4028 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_4027 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_4026 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_4025 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_4024 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_4023 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_4022 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_4021 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_4020 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_4019 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_4018 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_4017 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_4016 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_4015 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_4014 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_4013 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_4012 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_4011 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_4010 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_4009 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_4008 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4007 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_4006 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_4005 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_4004 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_4003 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV5 U1 ( .I(n2), .ZN(n3) );
  LVT_CLKNHSV4 U2 ( .I(n2), .ZN(n1) );
  LVT_CLKNHSV2 U3 ( .I(t_m_1_in), .ZN(n2) );
endmodule


module cell_2_128 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_4002 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4001 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4000 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3999 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3998 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3997 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3996 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3995 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3994 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3993 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3992 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3991 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3990 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3989 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3988 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3987 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3986 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3985 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3984 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3983 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3982 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3981 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3980 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3979 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3978 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3977 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3976 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3975 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n5), .A2(n6), .Z(t_i_out) );
endmodule


module cell_3_3974 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3973 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3972 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV4SR U1 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV4 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV2 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNHSV2P5 U5 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV4 U7 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_128 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_128 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_4002 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_4001 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_4000 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3999 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3998 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3997 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3996 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3995 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3994 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3993 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3992 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3991 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3990 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3989 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3988 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3987 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3986 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3985 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3984 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3983 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3982 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3981 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3980 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3979 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3978 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3977 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3976 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3975 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3974 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3973 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3972 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV3 U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV8SR U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_127 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3971 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3970 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3969 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3968 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3967 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3966 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3965 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3964 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3963 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3962 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3961 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3960 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3959 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_3958 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3957 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3956 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3955 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3954 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3953 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3952 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3951 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3950 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3949 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3948 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3947 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3946 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3945 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3944 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3943 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3942 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_3941 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV3SR U1 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV0SR U4 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U6 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U7 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_XNOR2HSV1 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_127 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1;

  cell_2_127 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_3971 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3970 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3969 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3968 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3967 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3966 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3965 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3964 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3963 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3962 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3961 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3960 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3959 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3958 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3957 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3956 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3955 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3954 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3953 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3952 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3951 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3950 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3949 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3948 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3947 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3946 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3945 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3944 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3943 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3942 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3941 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV2RT U1 ( .I(t_m_1_in), .Z(n1) );
endmodule


module cell_2_126 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_3940 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3939 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV1 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3938 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3937 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3936 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3935 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3934 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3933 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3932 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3931 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3930 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3929 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3928 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3927 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3926 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3925 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3924 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3923 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3922 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3921 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3920 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3919 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3918 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3917 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3916 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3915 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3914 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3913 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3912 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3911 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV2SR U5 ( .I(n10), .ZN(n4) );
  LVT_CLKNHSV0P5 U6 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV0P5 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_XOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
endmodule


module cell_3_3910 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2SR U4 ( .I(n9), .ZN(n2) );
  LVT_CLKNHSV0P5 U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV0P5 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV1 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_126 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_126 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3940 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3939 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3938 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3937 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3936 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3935 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3934 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3933 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3932 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3931 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3930 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3929 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3928 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3927 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3926 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3925 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3924 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3923 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3922 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3921 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3920 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3919 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3918 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3917 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3916 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3915 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3914 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3913 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3912 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3911 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3910 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV10 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV4SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_125 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3909 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3908 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3907 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3906 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3905 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3904 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3903 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3902 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3901 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3900 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3899 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3898 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3897 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3896 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3895 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3894 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3893 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3892 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3891 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3890 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3889 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3888 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3887 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3886 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3885 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3884 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3883 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3882 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3881 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_CLKNAND2HSV2 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV1 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNAND2HSV2 U3 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0SR U5 ( .I(n8), .ZN(n4) );
  LVT_INHSV2P5 U6 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV0 U7 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV2 U8 ( .A1(n10), .A2(n9), .Z(t_i_out) );
endmodule


module cell_3_3880 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_3879 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;

  LVT_INHSV2P5 U1 ( .I(n13), .ZN(n4) );
  LVT_NAND2HSV1 U2 ( .A1(n12), .A2(t_i_1_in), .ZN(n9) );
  LVT_INHSV0P5 U3 ( .I(t_i_1_in), .ZN(n8) );
  LVT_CLKNHSV2 U4 ( .I(n11), .ZN(n2) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  LVT_CLKNAND2HSV3 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n13) );
  LVT_NAND2HSV4 U7 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U8 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV1 U9 ( .A1(n7), .A2(n8), .ZN(n10) );
  LVT_NAND2HSV0P5 U10 ( .A1(n13), .A2(n11), .ZN(n5) );
  LVT_INHSV2 U11 ( .I(n12), .ZN(n7) );
  LVT_NAND2HSV0 U12 ( .A1(b_in), .A2(a_in), .ZN(n12) );
endmodule


module row_other_125 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_125 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_3909 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3908 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3907 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3906 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3905 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3904 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3903 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3902 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3901 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3900 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3899 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3898 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3897 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3896 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3895 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3894 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3893 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3892 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3891 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3890 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3889 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3888 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3887 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3886 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3885 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3884 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3883 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3882 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3881 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3880 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3879 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_124 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4, n5, n6, n7;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_INAND2HSV0 U1 ( .A1(n7), .B1(n6), .ZN(n5) );
  LVT_CLKNAND2HSV0 U2 ( .A1(n4), .A2(n5), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(n7), .A2(n3), .ZN(n4) );
  LVT_CLKNHSV0P5 U5 ( .I(n6), .ZN(n3) );
  LVT_CLKNAND2HSV1 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3878 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3877 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3876 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3875 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_OAI21HSV0 U2 ( .A1(n6), .A2(n4), .B(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(n6), .A2(n4), .ZN(n2) );
  LVT_XNOR2HSV1 U5 ( .A1(n5), .A2(t_i_1_in), .ZN(n4) );
endmodule


module cell_3_3874 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3873 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3872 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3871 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3870 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3869 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3868 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3867 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3866 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3865 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3864 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3863 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3862 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3861 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3860 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3859 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3858 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3857 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3856 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3855 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U4 ( .A1(n5), .A2(n2), .Z(t_i_out) );
endmodule


module cell_3_3854 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n8), .A2(n4), .ZN(n5) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(t_i_1_in), .ZN(n6) );
  LVT_NAND2HSV2 U4 ( .A1(n5), .A2(n6), .ZN(n7) );
  LVT_INHSV2 U5 ( .I(n8), .ZN(n2) );
  LVT_INHSV2 U6 ( .I(t_i_1_in), .ZN(n4) );
  LVT_XOR2HSV0 U7 ( .A1(n9), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
endmodule


module cell_3_3853 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3852 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3851 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n5), .A2(n2), .Z(t_i_out) );
endmodule


module cell_3_3850 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3849 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n2) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n5), .A2(n2), .Z(t_i_out) );
endmodule


module cell_3_3848 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_NAND2HSV2 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INAND2HSV2 U2 ( .A1(n9), .B1(n8), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n7), .A2(t_i_1_in), .Z(n8) );
  LVT_CLKNHSV0P5 U5 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0P5 U6 ( .A1(n9), .A2(n4), .ZN(n5) );
  LVT_NAND2HSV0P5 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
endmodule


module row_other_124 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_124 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_3878 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3877 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3876 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3875 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3874 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3873 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3872 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3871 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3870 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3869 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3868 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3867 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3866 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3865 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3864 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3863 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3862 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3861 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3860 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3859 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3858 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3857 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3856 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3855 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3854 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3853 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3852 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3851 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3850 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3849 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3848 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_4 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [31:0] a_in;
  input [31:0] g_in;
  input [31:0] b_in;
  input [31:0] t_m_1_in;
  input [30:0] t_i_1_in;
  input [30:0] t_i_2_in;
  output [31:0] a_out;
  output [31:0] g_out;
  output [30:0] t_i_1_out;
  output [30:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;
  wire   n1, n2, n4, n5, n7, n8, n10, n11, n13, n14, n16, n17, n19, n20, n22,
         n24, n25, n27, n29, n30, n31, n32, n33;
  wire   [30:0] t0;
  wire   [30:0] t1;
  wire   [30:0] t2;
  wire   [30:0] t3;
  wire   [30:0] t4;
  wire   [30:0] t5;
  wire   [30:0] t6;
  wire   [30:0] t7;
  wire   [30:0] t8;
  wire   [30:0] t9;
  wire   [30:0] t10;
  wire   [30:0] t11;
  wire   [30:0] t12;
  wire   [30:0] t13;
  wire   [30:0] t14;
  wire   [30:0] t15;
  wire   [30:0] t16;
  wire   [30:0] t17;
  wire   [30:0] t18;
  wire   [30:0] t19;
  wire   [30:0] t20;
  wire   [30:0] t21;
  wire   [30:0] t22;
  wire   [30:0] t23;
  wire   [30:0] t24;
  wire   [30:0] t25;
  wire   [30:0] t26;
  wire   [30:0] t27;
  wire   [30:0] t28;
  wire   [30:0] t29;
  wire   [30:0] t30;
  assign a_out[31] = a_in[31];
  assign a_out[30] = a_in[30];
  assign a_out[29] = a_in[29];
  assign a_out[28] = a_in[28];
  assign a_out[25] = a_in[25];
  assign a_out[23] = a_in[23];
  assign a_out[21] = a_in[21];
  assign a_out[20] = a_in[20];
  assign a_out[19] = a_in[19];
  assign a_out[18] = a_in[18];
  assign a_out[17] = a_in[17];
  assign a_out[16] = a_in[16];
  assign a_out[15] = a_in[15];
  assign a_out[14] = a_in[14];
  assign a_out[13] = a_in[13];
  assign a_out[12] = a_in[12];
  assign a_out[11] = a_in[11];
  assign a_out[10] = a_in[10];
  assign a_out[9] = a_in[9];
  assign a_out[8] = a_in[8];
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[30] = g_in[30];
  assign g_out[29] = g_in[29];
  assign g_out[27] = g_in[27];
  assign g_out[21] = g_in[21];
  assign g_out[20] = g_in[20];
  assign g_out[19] = g_in[19];
  assign g_out[18] = g_in[18];
  assign g_out[17] = g_in[17];
  assign g_out[16] = g_in[16];
  assign g_out[15] = g_in[15];
  assign g_out[14] = g_in[14];
  assign g_out[13] = g_in[13];
  assign g_out[12] = g_in[12];
  assign g_out[11] = g_in[11];
  assign g_out[10] = g_in[10];
  assign g_out[9] = g_in[9];
  assign g_out[8] = g_in[8];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_4 u0 ( .a_in({a_in[31:28], n20, n25, a_in[25], n8, a_in[23], n17, 
        a_in[21:0]}), .g_in({g_in[31:26], n14, n11, n2, n5, g_in[21:0]}), 
        .b_in(b_in[31]), .t_m_1_in(t_m_1_in[31]), .t_i_1_in({t_i_1_in, 
        t_i_1_in_0}), .t_i_2_in(t_i_2_in), .t_i_1_out(t0), .t_i_2_out(
        t_i_2_out[30]) );
  row_other_154 u1 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_in[31:29], g_out[28], 
        g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[30]), .t_m_1_in(
        t_m_1_in[30]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[29]) );
  row_other_153 u2 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_in[31:29], g_out[28], 
        g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[29]), .t_m_1_in(
        t_m_1_in[29]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[28]) );
  row_other_152 u3 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_in[31:29], g_out[28], 
        g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[28]), .t_m_1_in(
        t_m_1_in[28]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[27]) );
  row_other_151 u4 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[27]), 
        .t_m_1_in(t_m_1_in[27]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(
        t_i_2_out[26]) );
  row_other_150 u5 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[26]), 
        .t_m_1_in(t_m_1_in[26]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(
        t_i_2_out[25]) );
  row_other_149 u6 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[25]), 
        .t_m_1_in(t_m_1_in[25]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(
        t_i_2_out[24]) );
  row_other_148 u7 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[24]), 
        .t_m_1_in(t_m_1_in[24]), .t_i_1_in(t6), .t_i_1_out(t7), .t_i_2_out(
        t_i_2_out[23]) );
  row_other_147 u8 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[23]), 
        .t_m_1_in(n32), .t_i_1_in(t7), .t_i_1_out(t8), .t_i_2_out(
        t_i_2_out[22]) );
  row_other_146 u9 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[22]), 
        .t_m_1_in(t_m_1_in[22]), .t_i_1_in(t8), .t_i_1_out(t9), .t_i_2_out(
        t_i_2_out[21]) );
  row_other_145 u10 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[21]), 
        .t_m_1_in(t_m_1_in[21]), .t_i_1_in(t9), .t_i_1_out(t10), .t_i_2_out(
        t_i_2_out[20]) );
  row_other_144 u11 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[20]), 
        .t_m_1_in(t_m_1_in[20]), .t_i_1_in(t10), .t_i_1_out(t11), .t_i_2_out(
        t_i_2_out[19]) );
  row_other_143 u12 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[19]), 
        .t_m_1_in(t_m_1_in[19]), .t_i_1_in(t11), .t_i_1_out(t12), .t_i_2_out(
        t_i_2_out[18]) );
  row_other_142 u13 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[18]), 
        .t_m_1_in(t_m_1_in[18]), .t_i_1_in(t12), .t_i_1_out(t13), .t_i_2_out(
        t_i_2_out[17]) );
  row_other_141 u14 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[17]), 
        .t_m_1_in(t_m_1_in[17]), .t_i_1_in(t13), .t_i_1_out(t14), .t_i_2_out(
        t_i_2_out[16]) );
  row_other_140 u15 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[16]), 
        .t_m_1_in(t_m_1_in[16]), .t_i_1_in(t14), .t_i_1_out(t15), .t_i_2_out(
        t_i_2_out[15]) );
  row_other_139 u16 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[15]), 
        .t_m_1_in(t_m_1_in[15]), .t_i_1_in(t15), .t_i_1_out(t16), .t_i_2_out(
        t_i_2_out[14]) );
  row_other_138 u17 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[14]), 
        .t_m_1_in(t_m_1_in[14]), .t_i_1_in(t16), .t_i_1_out(t17), .t_i_2_out(
        t_i_2_out[13]) );
  row_other_137 u18 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[13]), 
        .t_m_1_in(t_m_1_in[13]), .t_i_1_in(t17), .t_i_1_out(t18), .t_i_2_out(
        t_i_2_out[12]) );
  row_other_136 u19 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[12]), 
        .t_m_1_in(t_m_1_in[12]), .t_i_1_in(t18), .t_i_1_out(t19), .t_i_2_out(
        t_i_2_out[11]) );
  row_other_135 u20 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[11]), 
        .t_m_1_in(t_m_1_in[11]), .t_i_1_in(t19), .t_i_1_out(t20), .t_i_2_out(
        t_i_2_out[10]) );
  row_other_134 u21 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[10]), 
        .t_m_1_in(n30), .t_i_1_in(t20), .t_i_1_out(t21), .t_i_2_out(
        t_i_2_out[9]) );
  row_other_133 u22 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[9]), 
        .t_m_1_in(t_m_1_in[9]), .t_i_1_in(t21), .t_i_1_out(t22), .t_i_2_out(
        t_i_2_out[8]) );
  row_other_132 u23 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[8]), 
        .t_m_1_in(t_m_1_in[8]), .t_i_1_in(t22), .t_i_1_out(t23), .t_i_2_out(
        t_i_2_out[7]) );
  row_other_131 u24 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[7]), 
        .t_m_1_in(t_m_1_in[7]), .t_i_1_in(t23), .t_i_1_out(t24), .t_i_2_out(
        t_i_2_out[6]) );
  row_other_130 u25 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[6]), 
        .t_m_1_in(t_m_1_in[6]), .t_i_1_in(t24), .t_i_1_out(t25), .t_i_2_out(
        t_i_2_out[5]) );
  row_other_129 u26 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[5]), 
        .t_m_1_in(t_m_1_in[5]), .t_i_1_in(t25), .t_i_1_out(t26), .t_i_2_out(
        t_i_2_out[4]) );
  row_other_128 u27 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[4]), 
        .t_m_1_in(t_m_1_in[4]), .t_i_1_in(t26), .t_i_1_out(t27), .t_i_2_out(
        t_i_2_out[3]) );
  row_other_127 u28 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[3]), 
        .t_m_1_in(t_m_1_in[3]), .t_i_1_in(t27), .t_i_1_out(t28), .t_i_2_out(
        t_i_2_out[2]) );
  row_other_126 u29 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[2]), 
        .t_m_1_in(t_m_1_in[2]), .t_i_1_in(t28), .t_i_1_out(t29), .t_i_2_out(
        t_i_2_out[1]) );
  row_other_125 u30 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[1]), 
        .t_m_1_in(t_m_1_in[1]), .t_i_1_in(t29), .t_i_1_out(t30), .t_i_2_out(
        t_i_2_out[0]) );
  row_other_124 u31 ( .a_in({a_in[31:28], a_out[27:26], a_in[25], a_out[24], 
        a_in[23], a_out[22], a_in[21:0]}), .g_in({g_out[31], g_in[30:29], 
        g_out[28], g_in[27], g_out[26:22], g_in[21:0]}), .b_in(b_in[0]), 
        .t_m_1_in(t_m_1_in[0]), .t_i_1_in(t30), .t_i_1_out(t_i_1_out), 
        .t_i_2_out(t_i_1_out_0) );
  LVT_INHSV10 U1 ( .I(n29), .ZN(n30) );
  LVT_INHSV2 U2 ( .I(n16), .ZN(n17) );
  LVT_INHSV2 U3 ( .I(n7), .ZN(n8) );
  LVT_INHSV2 U4 ( .I(a_in[22]), .ZN(n16) );
  LVT_INHSV2 U5 ( .I(a_in[24]), .ZN(n7) );
  LVT_INHSV2 U6 ( .I(a_in[27]), .ZN(n19) );
  LVT_INHSV2 U7 ( .I(g_in[22]), .ZN(n4) );
  LVT_INHSV2 U8 ( .I(g_in[23]), .ZN(n1) );
  LVT_INHSV2 U9 ( .I(g_in[24]), .ZN(n10) );
  LVT_INHSV2 U10 ( .I(g_in[25]), .ZN(n13) );
  LVT_CLKNHSV2 U11 ( .I(n1), .ZN(n2) );
  LVT_INHSV2SR U12 ( .I(n1), .ZN(g_out[23]) );
  LVT_INHSV2SR U13 ( .I(n4), .ZN(n5) );
  LVT_INHSV2SR U14 ( .I(n4), .ZN(g_out[22]) );
  LVT_INHSV2SR U15 ( .I(n7), .ZN(a_out[24]) );
  LVT_INHSV2SR U16 ( .I(n10), .ZN(n11) );
  LVT_INHSV2SR U17 ( .I(n10), .ZN(g_out[24]) );
  LVT_INHSV2SR U18 ( .I(n13), .ZN(n14) );
  LVT_INHSV2SR U19 ( .I(n13), .ZN(g_out[25]) );
  LVT_INHSV2SR U20 ( .I(n16), .ZN(a_out[22]) );
  LVT_INHSV2SR U21 ( .I(n19), .ZN(n20) );
  LVT_INHSV2SR U22 ( .I(n19), .ZN(a_out[27]) );
  LVT_INHSV8SR U23 ( .I(n31), .ZN(n32) );
  LVT_INHSV4 U24 ( .I(t_m_1_in[23]), .ZN(n31) );
  LVT_INHSV2 U25 ( .I(a_in[26]), .ZN(n24) );
  LVT_INHSV2 U26 ( .I(g_in[26]), .ZN(n22) );
  LVT_INHSV2 U27 ( .I(g_in[28]), .ZN(n27) );
  LVT_INHSV4SR U28 ( .I(t_m_1_in[10]), .ZN(n29) );
  LVT_INHSV2SR U29 ( .I(n22), .ZN(g_out[26]) );
  LVT_INHSV2SR U30 ( .I(n24), .ZN(n25) );
  LVT_INHSV2SR U31 ( .I(n24), .ZN(a_out[26]) );
  LVT_INHSV2SR U32 ( .I(n27), .ZN(g_out[28]) );
  LVT_CLKNHSV4 U33 ( .I(n33), .ZN(g_out[31]) );
  LVT_INHSV0SR U34 ( .I(g_in[31]), .ZN(n33) );
endmodule


module regist_32bit_25 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_32bit_24 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_31bit_16 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n1), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n2), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module PE_4 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro );
  input [31:0] a_in;
  input [31:0] g_in;
  input [31:0] b_in;
  input [30:0] t_i_1_in;
  input [30:0] t_i_2_in;
  output [31:0] a_out;
  output [31:0] g_out;
  output [31:0] b_out;
  output [30:0] t_i_1_out;
  output [30:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   n82, l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n74, n75, n76, n77, n78, n79, n80, n81;
  wire   [31:0] l_a;
  wire   [31:0] l_g;
  wire   [30:0] l_t_i_1_in;
  wire   [30:0] l_t_i_2_in;
  wire   [31:0] mux_b;
  wire   [31:0] mux_bq;
  wire   [30:0] to_7;
  wire   [30:0] ti_7;
  wire   [31:0] ao;
  wire   [31:0] go;
  wire   [30:0] to;

  LVT_AO22HSV0 U39 ( .A1(mux_bq[5]), .A2(n69), .B1(b_out[5]), .B2(n35), .Z(
        mux_b[5]) );
  LVT_AO22HSV0 U40 ( .A1(mux_bq[4]), .A2(n69), .B1(b_out[4]), .B2(n35), .Z(
        mux_b[4]) );
  LVT_AO22HSV0 U41 ( .A1(mux_bq[3]), .A2(n69), .B1(b_out[3]), .B2(n35), .Z(
        mux_b[3]) );
  LVT_AO22HSV0 U44 ( .A1(mux_bq[2]), .A2(n69), .B1(b_out[2]), .B2(n35), .Z(
        mux_b[2]) );
  LVT_AO22HSV0 U55 ( .A1(mux_bq[1]), .A2(n69), .B1(b_out[1]), .B2(n35), .Z(
        mux_b[1]) );
  LVT_AO22HSV0 U64 ( .A1(mux_bq[11]), .A2(n69), .B1(b_out[11]), .B2(n35), .Z(
        mux_b[11]) );
  LVT_AO22HSV0 U65 ( .A1(mux_bq[10]), .A2(n69), .B1(b_out[10]), .B2(n35), .Z(
        mux_b[10]) );
  LVT_AO22HSV0 U66 ( .A1(mux_bq[0]), .A2(n69), .B1(b_out[0]), .B2(n35), .Z(
        mux_b[0]) );
  LVT_NOR2HSV0 U67 ( .A1(n2), .A2(n3), .ZN(c_t_i_1_in_0) );
  LVT_AOI21HSV0 U69 ( .A1(n4), .A2(n5), .B(n3), .ZN(\c_t_i_1_in[0] ) );
  LVT_AND4HSV0 U71 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .Z(n5) );
  LVT_NOR4HSV0 U72 ( .A1(l_t_i_1_in[9]), .A2(l_t_i_1_in[8]), .A3(l_t_i_1_in[7]), .A4(l_t_i_1_in[6]), .ZN(n9) );
  LVT_NOR4HSV0 U73 ( .A1(l_t_i_1_in[5]), .A2(l_t_i_1_in[4]), .A3(l_t_i_1_in[3]), .A4(l_t_i_1_in[30]), .ZN(n8) );
  LVT_NOR4HSV0 U74 ( .A1(l_t_i_1_in[2]), .A2(l_t_i_1_in[29]), .A3(
        l_t_i_1_in[28]), .A4(l_t_i_1_in[27]), .ZN(n7) );
  LVT_NOR4HSV0 U75 ( .A1(l_t_i_1_in[26]), .A2(l_t_i_1_in[25]), .A3(
        l_t_i_1_in[24]), .A4(l_t_i_1_in[23]), .ZN(n6) );
  LVT_AND4HSV0 U76 ( .A1(n10), .A2(n11), .A3(n12), .A4(n13), .Z(n4) );
  LVT_NOR4HSV0 U77 ( .A1(l_t_i_1_in[22]), .A2(l_t_i_1_in[21]), .A3(
        l_t_i_1_in[20]), .A4(l_t_i_1_in[1]), .ZN(n13) );
  LVT_NOR4HSV0 U78 ( .A1(l_t_i_1_in[19]), .A2(l_t_i_1_in[18]), .A3(
        l_t_i_1_in[17]), .A4(l_t_i_1_in[16]), .ZN(n12) );
  LVT_NOR4HSV0 U79 ( .A1(l_t_i_1_in[15]), .A2(l_t_i_1_in[14]), .A3(
        l_t_i_1_in[13]), .A4(l_t_i_1_in[12]), .ZN(n11) );
  LVT_NOR3HSV0 U80 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[11]), .A3(
        l_t_i_1_in[10]), .ZN(n10) );
  regist_32bit_29 u0 ( .clk(clk), .rstn(n80), .in(a_in), .out(l_a) );
  regist_32bit_28 u1 ( .clk(clk), .rstn(n80), .in(b_in), .out(b_out) );
  regist_32bit_27 u2 ( .clk(clk), .rstn(n80), .in(g_in), .out(l_g) );
  regist_1bit_19 u3 ( .clk(clk), .rstn(n80), .in(ctr), .out(l_ctr) );
  regist_1bit_18 u4 ( .clk(clk), .rstn(n80), .in(n69), .out(ctro) );
  regist_31bit_19 u5 ( .clk(clk), .rstn(n80), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_31bit_18 u6 ( .clk(clk), .rstn(n80), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_17 u7 ( .clk(clk), .rstn(n80), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_32bit_26 u9 ( .clk(clk), .rstn(n80), .in(mux_b), .out(mux_bq) );
  regist_1bit_16 u10 ( .clk(clk), .rstn(n80), .in(to_1), .out(ti_1) );
  regist_31bit_17 u11 ( .clk(clk), .rstn(n80), .in({to_7[30], n74, to_7[28:25], 
        n39, to_7[23:14], n20, to_7[12:5], n71, to_7[3:0]}), .out(ti_7) );
  PE_core_4 pe ( .a_in({l_a[31:30], n22, l_a[28:0]}), .g_in(l_g), .b_in(mux_bq), .t_m_1_in({to_1, to_7[30], n74, to_7[28:25], n39, to_7[23:5], n71, to_7[3:0]}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out({t_i_2_out[30:12], n82, 
        t_i_2_out[10:0]}), .t_i_1_out_0(t_i_1_out_0) );
  regist_32bit_25 u12 ( .clk(clk), .rstn(n80), .in(ao), .out(a_out) );
  regist_32bit_24 u13 ( .clk(clk), .rstn(n80), .in(go), .out(g_out) );
  regist_31bit_16 u14 ( .clk(clk), .rstn(n80), .in(to), .out(t_i_1_out) );
  LVT_OR2HSV16RD U2 ( .A1(n45), .A2(n44), .Z(to_7[9]) );
  LVT_CLKNHSV12 U3 ( .I(l_ctr), .ZN(n79) );
  LVT_CLKNHSV8 U4 ( .I(n14), .ZN(to_7[21]) );
  LVT_CLKNAND2HSV3 U5 ( .A1(t_i_2_out[7]), .A2(n18), .ZN(n43) );
  LVT_NAND2HSV4 U6 ( .A1(n65), .A2(n64), .ZN(to_7[12]) );
  LVT_NAND2HSV8 U7 ( .A1(n42), .A2(n43), .ZN(to_7[7]) );
  LVT_CLKNAND2HSV2 U8 ( .A1(t_i_2_out[22]), .A2(n18), .ZN(n55) );
  LVT_INHSV6SR U9 ( .I(n66), .ZN(n74) );
  LVT_NAND2HSV12 U10 ( .A1(n29), .A2(n30), .ZN(to_7[13]) );
  LVT_CLKNAND2HSV3 U11 ( .A1(t_i_2_out[20]), .A2(n18), .ZN(n16) );
  LVT_NOR2HSV8 U12 ( .A1(n46), .A2(n47), .ZN(n14) );
  LVT_BUFHSV4 U13 ( .I(n1), .Z(n18) );
  LVT_INHSV2 U14 ( .I(ctro), .ZN(n1) );
  LVT_NAND2HSV2 U15 ( .A1(ti_7[10]), .A2(ctro), .ZN(n23) );
  LVT_NAND2HSV4 U16 ( .A1(n76), .A2(n75), .ZN(to_7[16]) );
  LVT_CLKNAND2HSV4 U17 ( .A1(n61), .A2(n60), .ZN(to_7[11]) );
  LVT_CLKNAND2HSV3 U18 ( .A1(n82), .A2(n18), .ZN(n61) );
  LVT_NAND2HSV4 U19 ( .A1(ti_7[20]), .A2(ctro), .ZN(n15) );
  LVT_NAND2HSV4 U20 ( .A1(n15), .A2(n16), .ZN(to_7[20]) );
  LVT_CLKNAND2HSV8 U21 ( .A1(n36), .A2(n37), .ZN(to_7[0]) );
  LVT_AND2HSV8 U22 ( .A1(t_i_2_out[30]), .A2(n17), .Z(n68) );
  LVT_CLKBUFHSV5 U23 ( .I(n1), .Z(n17) );
  LVT_NAND2HSV2 U24 ( .A1(t_i_2_out[6]), .A2(n18), .ZN(n51) );
  LVT_CLKNHSV4 U25 ( .I(n21), .ZN(n22) );
  LVT_INHSV2 U26 ( .I(l_a[29]), .ZN(n21) );
  LVT_CLKNAND2HSV8 U27 ( .A1(n32), .A2(n31), .ZN(to_7[3]) );
  LVT_NAND2HSV2 U28 ( .A1(ti_7[23]), .A2(ctro), .ZN(n25) );
  LVT_INHSV4 U29 ( .I(n38), .ZN(n39) );
  LVT_INHSV0SR U30 ( .I(to_7[13]), .ZN(n19) );
  LVT_INHSV2 U31 ( .I(n19), .ZN(n20) );
  LVT_AO22HSV2 U32 ( .A1(mux_bq[15]), .A2(l_ctr), .B1(b_out[15]), .B2(n3), .Z(
        mux_b[15]) );
  LVT_AO22HSV2 U33 ( .A1(mux_bq[25]), .A2(l_ctr), .B1(b_out[25]), .B2(n35), 
        .Z(mux_b[25]) );
  LVT_AO22HSV2 U34 ( .A1(mux_bq[12]), .A2(l_ctr), .B1(b_out[12]), .B2(n3), .Z(
        mux_b[12]) );
  LVT_AO22HSV2 U35 ( .A1(mux_bq[13]), .A2(l_ctr), .B1(b_out[13]), .B2(n3), .Z(
        mux_b[13]) );
  LVT_AO22HSV2 U36 ( .A1(mux_bq[14]), .A2(l_ctr), .B1(b_out[14]), .B2(n3), .Z(
        mux_b[14]) );
  LVT_AO22HSV2 U37 ( .A1(mux_bq[17]), .A2(l_ctr), .B1(b_out[17]), .B2(n3), .Z(
        mux_b[17]) );
  LVT_AO22HSV2 U38 ( .A1(mux_bq[18]), .A2(l_ctr), .B1(b_out[18]), .B2(n3), .Z(
        mux_b[18]) );
  LVT_AO22HSV2 U42 ( .A1(mux_bq[19]), .A2(l_ctr), .B1(b_out[19]), .B2(n3), .Z(
        mux_b[19]) );
  LVT_AO22HSV2 U43 ( .A1(mux_bq[20]), .A2(l_ctr), .B1(b_out[20]), .B2(n3), .Z(
        mux_b[20]) );
  LVT_AO22HSV2 U45 ( .A1(mux_bq[21]), .A2(l_ctr), .B1(b_out[21]), .B2(n3), .Z(
        mux_b[21]) );
  LVT_AO22HSV2 U46 ( .A1(mux_bq[22]), .A2(l_ctr), .B1(b_out[22]), .B2(n3), .Z(
        mux_b[22]) );
  LVT_AO22HSV2 U47 ( .A1(mux_bq[23]), .A2(l_ctr), .B1(b_out[23]), .B2(n35), 
        .Z(mux_b[23]) );
  LVT_AO22HSV2 U48 ( .A1(mux_bq[26]), .A2(l_ctr), .B1(b_out[26]), .B2(n35), 
        .Z(mux_b[26]) );
  LVT_AO22HSV2 U49 ( .A1(mux_bq[28]), .A2(l_ctr), .B1(b_out[28]), .B2(n3), .Z(
        mux_b[28]) );
  LVT_AO22HSV2 U50 ( .A1(mux_bq[30]), .A2(l_ctr), .B1(b_out[30]), .B2(n3), .Z(
        mux_b[30]) );
  LVT_AO22HSV2 U51 ( .A1(mux_bq[6]), .A2(l_ctr), .B1(b_out[6]), .B2(n35), .Z(
        mux_b[6]) );
  LVT_AO22HSV2 U52 ( .A1(mux_bq[7]), .A2(l_ctr), .B1(b_out[7]), .B2(n35), .Z(
        mux_b[7]) );
  LVT_AO22HSV2 U53 ( .A1(mux_bq[8]), .A2(l_ctr), .B1(b_out[8]), .B2(n35), .Z(
        mux_b[8]) );
  LVT_AO22HSV2 U54 ( .A1(mux_bq[9]), .A2(l_ctr), .B1(b_out[9]), .B2(n35), .Z(
        mux_b[9]) );
  LVT_AO22HSV2 U56 ( .A1(mux_bq[16]), .A2(l_ctr), .B1(b_out[16]), .B2(n3), .Z(
        mux_b[16]) );
  LVT_AO22HSV2 U57 ( .A1(mux_bq[24]), .A2(l_ctr), .B1(b_out[24]), .B2(n35), 
        .Z(mux_b[24]) );
  LVT_AO22HSV2 U58 ( .A1(mux_bq[27]), .A2(l_ctr), .B1(b_out[27]), .B2(n35), 
        .Z(mux_b[27]) );
  LVT_AO22HSV2 U59 ( .A1(mux_bq[29]), .A2(l_ctr), .B1(b_out[29]), .B2(n3), .Z(
        mux_b[29]) );
  LVT_OR2HSV12RD U60 ( .A1(n59), .A2(n58), .Z(to_7[5]) );
  LVT_CLKNAND2HSV3 U61 ( .A1(n23), .A2(n24), .ZN(to_7[10]) );
  LVT_OR2HSV12RD U62 ( .A1(n48), .A2(n49), .Z(to_7[14]) );
  LVT_NAND2HSV4 U63 ( .A1(t_i_2_out[17]), .A2(n18), .ZN(n57) );
  LVT_CLKAND2HSV4 U68 ( .A1(t_i_2_out[5]), .A2(n18), .Z(n59) );
  LVT_CLKAND2HSV4 U70 ( .A1(t_i_2_out[14]), .A2(n18), .Z(n49) );
  LVT_NAND2HSV4 U81 ( .A1(t_i_2_out[16]), .A2(n18), .ZN(n76) );
  LVT_CLKNAND2HSV3 U82 ( .A1(t_i_2_out[12]), .A2(n18), .ZN(n65) );
  LVT_CLKNAND2HSV3 U83 ( .A1(t_i_2_out[27]), .A2(n18), .ZN(n41) );
  LVT_CLKNAND2HSV8 U84 ( .A1(n56), .A2(n57), .ZN(to_7[17]) );
  LVT_NAND2HSV4 U85 ( .A1(t_i_2_out[23]), .A2(n18), .ZN(n26) );
  LVT_NAND2HSV4 U86 ( .A1(n52), .A2(n53), .ZN(to_7[26]) );
  LVT_CLKNAND2HSV3 U87 ( .A1(t_i_2_out[26]), .A2(n18), .ZN(n53) );
  LVT_CLKNAND2HSV3 U88 ( .A1(t_i_2_out[10]), .A2(n18), .ZN(n24) );
  LVT_NAND2HSV4 U89 ( .A1(t_i_2_out[3]), .A2(n18), .ZN(n32) );
  LVT_NAND2HSV4 U90 ( .A1(n25), .A2(n26), .ZN(to_7[23]) );
  LVT_CLKNAND2HSV2 U91 ( .A1(ti_7[2]), .A2(ctro), .ZN(n27) );
  LVT_CLKNAND2HSV3 U92 ( .A1(t_i_2_out[2]), .A2(n18), .ZN(n28) );
  LVT_NAND2HSV4 U93 ( .A1(n27), .A2(n28), .ZN(to_7[2]) );
  LVT_CLKNAND2HSV4 U94 ( .A1(n41), .A2(n40), .ZN(to_7[27]) );
  LVT_CLKNAND2HSV8 U95 ( .A1(n34), .A2(n33), .ZN(to_7[8]) );
  LVT_CLKNAND2HSV4 U96 ( .A1(n54), .A2(n55), .ZN(to_7[22]) );
  LVT_AO22HSV2 U97 ( .A1(mux_bq[31]), .A2(l_ctr), .B1(b_out[31]), .B2(n3), .Z(
        mux_b[31]) );
  LVT_NAND2HSV8 U98 ( .A1(t_i_2_out[13]), .A2(n18), .ZN(n30) );
  LVT_NAND2HSV4 U99 ( .A1(t_i_2_out[8]), .A2(n18), .ZN(n34) );
  LVT_INHSV2 U100 ( .I(n81), .ZN(n80) );
  LVT_NAND2HSV2 U101 ( .A1(ti_7[13]), .A2(ctro), .ZN(n29) );
  LVT_NAND2HSV2 U102 ( .A1(ti_7[3]), .A2(ctro), .ZN(n31) );
  LVT_NAND2HSV2 U103 ( .A1(ti_7[8]), .A2(ctro), .ZN(n33) );
  LVT_NAND2HSV4 U104 ( .A1(n51), .A2(n50), .ZN(to_7[6]) );
  LVT_INHSV2 U105 ( .I(n69), .ZN(n35) );
  LVT_CLKNAND2HSV8 U106 ( .A1(n77), .A2(n78), .ZN(to_1) );
  LVT_INHSV4 U107 ( .I(n70), .ZN(n71) );
  LVT_NAND2HSV0 U108 ( .A1(ti_7[0]), .A2(ctro), .ZN(n36) );
  LVT_CLKNAND2HSV4 U109 ( .A1(t_i_2_out[0]), .A2(n18), .ZN(n37) );
  LVT_NAND2HSV4 U110 ( .A1(ti_1), .A2(l_ctr), .ZN(n77) );
  LVT_CLKNAND2HSV8 U111 ( .A1(n79), .A2(l_t_i_1_in_0), .ZN(n78) );
  LVT_AOI22HSV4 U112 ( .A1(ti_7[24]), .A2(ctro), .B1(t_i_2_out[24]), .B2(n18), 
        .ZN(n38) );
  LVT_NAND2HSV0 U113 ( .A1(ti_7[27]), .A2(ctro), .ZN(n40) );
  LVT_NAND2HSV0 U114 ( .A1(ti_7[7]), .A2(ctro), .ZN(n42) );
  LVT_AND2HSV0RD U115 ( .A1(ti_7[9]), .A2(ctro), .Z(n44) );
  LVT_AND2HSV8 U116 ( .A1(t_i_2_out[9]), .A2(n18), .Z(n45) );
  LVT_AND2HSV0RD U117 ( .A1(ti_7[21]), .A2(ctro), .Z(n46) );
  LVT_AND2HSV8 U118 ( .A1(t_i_2_out[21]), .A2(n18), .Z(n47) );
  LVT_AND2HSV0RD U119 ( .A1(ti_7[14]), .A2(ctro), .Z(n48) );
  LVT_NAND2HSV0 U120 ( .A1(ti_7[6]), .A2(ctro), .ZN(n50) );
  LVT_INHSV0SR U121 ( .I(l_ctr), .ZN(n3) );
  LVT_NAND2HSV0 U122 ( .A1(ti_7[26]), .A2(ctro), .ZN(n52) );
  LVT_NAND2HSV0 U123 ( .A1(ti_7[22]), .A2(ctro), .ZN(n54) );
  LVT_NAND2HSV0 U124 ( .A1(ti_7[17]), .A2(ctro), .ZN(n56) );
  LVT_AND2HSV0RD U125 ( .A1(ti_7[5]), .A2(ctro), .Z(n58) );
  LVT_NAND2HSV0 U126 ( .A1(ti_7[11]), .A2(ctro), .ZN(n60) );
  LVT_AND2HSV0RD U127 ( .A1(ti_7[1]), .A2(ctro), .Z(n62) );
  LVT_AND2HSV8 U128 ( .A1(t_i_2_out[1]), .A2(n18), .Z(n63) );
  LVT_OR2HSV16RD U129 ( .A1(n63), .A2(n62), .Z(to_7[1]) );
  LVT_NAND2HSV0 U130 ( .A1(ti_7[12]), .A2(ctro), .ZN(n64) );
  LVT_AOI22HSV4 U131 ( .A1(ti_7[29]), .A2(ctro), .B1(t_i_2_out[29]), .B2(n18), 
        .ZN(n66) );
  LVT_AND2HSV0RD U132 ( .A1(ti_7[30]), .A2(ctro), .Z(n67) );
  LVT_OR2HSV16RD U133 ( .A1(n68), .A2(n67), .Z(to_7[30]) );
  LVT_BUFHSV2RT U134 ( .I(l_ctr), .Z(n69) );
  LVT_AOI22HSV4 U135 ( .A1(ti_7[4]), .A2(ctro), .B1(t_i_2_out[4]), .B2(n18), 
        .ZN(n70) );
  LVT_INHSV0SR U136 ( .I(n82), .ZN(n72) );
  LVT_INHSV2 U137 ( .I(n72), .ZN(t_i_2_out[11]) );
  LVT_AO22HSV4 U138 ( .A1(ti_7[15]), .A2(ctro), .B1(t_i_2_out[15]), .B2(n18), 
        .Z(to_7[15]) );
  LVT_NAND2HSV0 U139 ( .A1(ti_7[16]), .A2(ctro), .ZN(n75) );
  LVT_AO22HSV4 U140 ( .A1(ti_7[19]), .A2(ctro), .B1(t_i_2_out[19]), .B2(n18), 
        .Z(to_7[19]) );
  LVT_AO22HSV4 U141 ( .A1(ti_7[18]), .A2(ctro), .B1(t_i_2_out[18]), .B2(n18), 
        .Z(to_7[18]) );
  LVT_AO22HSV4 U142 ( .A1(ti_7[28]), .A2(ctro), .B1(t_i_2_out[28]), .B2(n18), 
        .Z(to_7[28]) );
  LVT_AO22HSV4 U143 ( .A1(ti_7[25]), .A2(ctro), .B1(t_i_2_out[25]), .B2(n18), 
        .Z(to_7[25]) );
  LVT_INHSV1 U144 ( .I(l_t_i_1_in_0), .ZN(n2) );
  LVT_INHSV2 U145 ( .I(rstn), .ZN(n81) );
endmodule


module regist_32bit_23 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV4 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n2), .Q(out[31]) );
  LVT_DRNQHSV4 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n2), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n1), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n1), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n1), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n1), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n1), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n1), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n1), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n2), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n2), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n2), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_CLKNHSV4 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_32bit_22 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV2 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n2), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n2), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n2), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_32bit_21 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n8, n9, n1, n3, n5, n6, n7;

  LVT_DRNQHSV4 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n5), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n6), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n5), .Q(n9) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n5), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n5), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n5), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n6), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n6), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n5), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n5), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n5), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n5), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n5), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n5), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n5), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n5), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n5), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n5), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n5), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n5), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n6), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n6), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n6), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n6), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n6), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n6), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n6), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n5), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n5), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n5), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n5), .Q(out[29]) );
  LVT_DRNQHSV4 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n6), .Q(n8) );
  LVT_CLKNHSV8 U3 ( .I(n8), .ZN(n3) );
  LVT_INHSV8SR U4 ( .I(n1), .ZN(out[30]) );
  LVT_INHSV24SR U5 ( .I(n3), .ZN(out[31]) );
  LVT_INHSV2 U6 ( .I(n9), .ZN(n1) );
  LVT_INHSV2 U7 ( .I(rstn), .ZN(n7) );
  LVT_INHSV2 U8 ( .I(n7), .ZN(n6) );
  LVT_CLKNHSV4 U9 ( .I(n7), .ZN(n5) );
endmodule


module regist_1bit_15 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_14 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_31bit_15 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n1), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n1), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n1), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n1), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n1), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n1), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n1), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n2) );
  LVT_CLKNHSV4 U4 ( .I(n2), .ZN(n1) );
endmodule


module regist_31bit_14 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n1), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(rstn), .Q(out[25])
         );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n1), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n1), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n1), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n1), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(rstn), .Q(out[24])
         );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n1), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n1), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n2) );
  LVT_CLKNHSV4 U4 ( .I(n2), .ZN(n1) );
endmodule


module regist_1bit_13 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_32bit_20 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n2), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n2), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n2), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n2), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n2), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n2), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n2), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_CLKNHSV4 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_1bit_12 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_31bit_13 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n2), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n2), .Q(out[28]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n2), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n2), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n2), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n2), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n1) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n2) );
endmodule


module cell_3_3847 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_123 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_122 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_121 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_120 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_119 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_118 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_117 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_116 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_115 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_114 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_113 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_112 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_111 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_110 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_109 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_108 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_107 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_106 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_105 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_104 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_103 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_102 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV1 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_101 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_100 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_99 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_98 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_XOR3HSV1 U2 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
endmodule


module cell_4_97 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_96 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_95 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
endmodule


module cell_4_94 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV2 U1 ( .A1(n5), .A2(n2), .A3(n4), .Z(t_i_out) );
  LVT_CLKNAND2HSV3 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_93 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n3, n5, n6, n7;

  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_OAI21HSV2 U2 ( .A1(n7), .A2(n5), .B(n2), .ZN(t_i_out) );
  LVT_NAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .ZN(n3) );
  LVT_NAND2HSV2 U4 ( .A1(n7), .A2(n5), .ZN(n2) );
  LVT_XNOR2HSV4 U6 ( .A1(n3), .A2(n6), .ZN(n5) );
endmodule


module row_1_3 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [31:0] t_i_1_in;
  input [30:0] t_i_2_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_3_3847 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_123 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(t_i_1_out[1])
         );
  cell_4_122 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(t_i_1_out[2])
         );
  cell_4_121 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(t_i_1_out[3])
         );
  cell_4_120 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(t_i_1_out[4])
         );
  cell_4_119 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(t_i_1_out[5])
         );
  cell_4_118 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(t_i_1_out[6])
         );
  cell_4_117 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(t_i_1_out[7])
         );
  cell_4_116 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_2_in(t_i_2_in[7]), .t_i_out(t_i_1_out[8])
         );
  cell_4_115 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[9]), .t_i_2_in(t_i_2_in[8]), .t_i_out(t_i_1_out[9])
         );
  cell_4_114 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[10]), .t_i_2_in(t_i_2_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_4_113 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[11]), .t_i_2_in(t_i_2_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_4_112 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[12]), .t_i_2_in(t_i_2_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_4_111 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[13]), .t_i_2_in(t_i_2_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_4_110 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[14]), .t_i_2_in(t_i_2_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_4_109 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[15]), .t_i_2_in(t_i_2_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_4_108 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[16]), .t_i_2_in(t_i_2_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_4_107 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[17]), .t_i_2_in(t_i_2_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_4_106 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[18]), .t_i_2_in(t_i_2_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_4_105 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[19]), .t_i_2_in(t_i_2_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_4_104 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[20]), .t_i_2_in(t_i_2_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_4_103 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[21]), .t_i_2_in(t_i_2_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_4_102 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[22]), .t_i_2_in(t_i_2_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_4_101 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[23]), .t_i_2_in(t_i_2_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_4_100 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_2_in(t_i_2_in[23]), .t_i_out(
        t_i_1_out[24]) );
  cell_4_99 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_2_in(t_i_2_in[24]), .t_i_out(
        t_i_1_out[25]) );
  cell_4_98 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[26]), .t_i_2_in(t_i_2_in[25]), .t_i_out(
        t_i_1_out[26]) );
  cell_4_97 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_2_in(t_i_2_in[26]), .t_i_out(
        t_i_1_out[27]) );
  cell_4_96 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_2_in(t_i_2_in[27]), .t_i_out(
        t_i_1_out[28]) );
  cell_4_95 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_2_in(t_i_2_in[28]), .t_i_out(
        t_i_1_out[29]) );
  cell_4_94 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_2_in(t_i_2_in[29]), .t_i_out(
        t_i_1_out[30]) );
  cell_4_93 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[31]), .t_i_2_in(t_i_2_in[30]), .t_i_out(
        t_i_2_out) );
  LVT_CLKNHSV6 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV2SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_123 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3846 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3845 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3844 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3843 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3842 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3841 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3840 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3839 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3838 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3837 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3836 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3835 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3834 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3833 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3832 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3831 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3830 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3829 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3828 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3827 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3826 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3825 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3824 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3823 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n5), .A2(n6), .Z(t_i_out) );
endmodule


module cell_3_3822 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3821 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3820 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3819 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV3 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3818 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0P5 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_CLKNHSV0P5 U5 ( .I(n10), .ZN(n4) );
  LVT_CLKNHSV2 U6 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV0 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_XOR2HSV2 U8 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
endmodule


module cell_3_3817 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3816 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_123 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_123 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3846 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3845 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3844 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3843 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3842 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3841 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3840 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3839 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3838 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3837 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3836 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3835 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3834 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3833 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3832 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3831 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3830 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3829 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3828 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3827 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3826 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3825 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3824 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3823 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3822 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3821 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3820 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3819 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3818 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3817 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3816 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2P5 U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV8 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_122 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3815 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3814 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3813 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3812 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3811 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3810 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3809 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3808 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3807 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3806 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3805 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3804 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3803 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3802 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3801 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3800 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3799 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3798 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3797 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3796 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3795 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3794 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3793 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3792 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3791 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3790 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3789 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3788 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3787 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3786 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV1 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module cell_3_3785 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n1, n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(t_i_1_in), .ZN(n4) );
  LVT_OAI21HSV2 U2 ( .A1(n1), .A2(n4), .B(n2), .ZN(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(n1), .A2(n4), .ZN(n2) );
  LVT_NAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n1) );
endmodule


module row_other_122 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_2_122 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3815 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3814 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3813 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3812 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3811 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3810 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3809 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3808 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3807 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3806 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3805 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3804 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3803 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3802 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3801 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3800 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3799 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3798 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3797 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3796 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3795 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3794 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3793 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3792 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3791 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3790 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3789 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3788 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3787 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3786 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3785 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV2P5 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV6 U2 ( .I(t_m_1_in), .ZN(n1) );
  LVT_CLKNHSV8 U3 ( .I(n1), .ZN(n3) );
  LVT_CLKNHSV3 U4 ( .I(n1), .ZN(n4) );
endmodule


module cell_2_121 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3784 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3783 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3782 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3781 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3780 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3779 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3778 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3777 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3776 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3775 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3774 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3773 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3772 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3771 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3770 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3769 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3768 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3767 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3766 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3765 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3764 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3763 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3762 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3761 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3760 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3759 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3758 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3757 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3756 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3755 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV2 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV1 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U3 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0SR U4 ( .I(n8), .ZN(n4) );
  LVT_CLKNHSV2P5 U5 ( .I(t_i_1_in), .ZN(n5) );
  LVT_CLKNAND2HSV8 U6 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV2 U7 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_3754 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_121 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_121 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_3784 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3783 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3782 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3781 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3780 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3779 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3778 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3777 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3776 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3775 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3774 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3773 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3772 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3771 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3770 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3769 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3768 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3767 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3766 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3765 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3764 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3763 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3762 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3761 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3760 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3759 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3758 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3757 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3756 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3755 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3754 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_120 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_3753 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3752 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3751 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3750 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3749 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3748 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3747 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3746 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3745 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3744 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3743 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3742 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3741 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3740 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3739 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3738 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3737 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3736 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3735 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3734 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3733 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3732 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3731 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3730 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3729 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV0P5 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U3 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0SR U5 ( .I(n8), .ZN(n4) );
  LVT_CLKNHSV2 U6 ( .I(t_i_1_in), .ZN(n5) );
  LVT_CLKNAND2HSV4 U7 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV2 U8 ( .A1(n10), .A2(n9), .Z(t_i_out) );
endmodule


module cell_3_3728 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3727 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3726 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3725 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKXOR2HSV2 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3724 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0P5 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_CLKNHSV0P5 U5 ( .I(n10), .ZN(n4) );
  LVT_INHSV0P5 U6 ( .I(n9), .ZN(n5) );
  LVT_XOR2HSV2 U7 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_NAND2HSV0 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_3723 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV4 U2 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV0P5 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNHSV2 U7 ( .I(n9), .ZN(n2) );
  LVT_INHSV2 U8 ( .I(n7), .ZN(n4) );
endmodule


module row_other_120 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_120 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3753 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3752 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3751 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3750 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3749 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3748 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3747 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3746 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3745 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3744 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3743 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3742 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3741 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3740 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3739 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3738 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3737 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3736 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3735 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3734 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3733 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3732 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3731 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3730 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3729 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3728 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3727 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3726 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3725 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3724 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3723 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV4 U1 ( .I(n1), .ZN(n2) );
  LVT_CLKNHSV1 U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_119 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_3722 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3721 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3720 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3719 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3718 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3717 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3716 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3715 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3714 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3713 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3712 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3711 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3710 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3709 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3708 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3707 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3706 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3705 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3704 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3703 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3702 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3701 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3700 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3699 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3698 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3697 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3696 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV1 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U3 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_CLKNHSV0P5 U4 ( .I(n8), .ZN(n4) );
  LVT_INHSV2 U5 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV4 U6 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV2 U7 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_3695 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3694 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U3 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_CLKNAND2HSV1 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U5 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_3_3693 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3692 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_OAI21HSV2 U2 ( .A1(n6), .A2(n4), .B(n2), .ZN(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(n6), .A2(n4), .ZN(n2) );
  LVT_XNOR2HSV4 U5 ( .A1(n5), .A2(t_i_1_in), .ZN(n4) );
endmodule


module row_other_119 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_119 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3722 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3721 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3720 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3719 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3718 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3717 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3716 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3715 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3714 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3713 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3712 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3711 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3710 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3709 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3708 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3707 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3706 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3705 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3704 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3703 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3702 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3701 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3700 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3699 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3698 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3697 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3696 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3695 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3694 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3693 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3692 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV2 U1 ( .I(t_m_1_in), .ZN(n2) );
  LVT_INHSV6 U2 ( .I(n2), .ZN(n1) );
endmodule


module cell_2_118 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3691 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3690 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3689 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3688 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3687 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3686 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3685 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3684 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3683 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3682 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3681 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3680 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3679 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3678 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3677 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3676 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3675 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3674 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3673 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3672 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3671 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3670 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3669 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3668 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3667 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3666 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3665 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3664 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3663 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV2 U1 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0P5 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_CLKNHSV0 U5 ( .I(n10), .ZN(n4) );
  LVT_INHSV2P5 U6 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV0P5 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_XOR2HSV2 U8 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
endmodule


module cell_3_3662 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3661 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNHSV0P5 U2 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV0 U5 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2SR U6 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV2 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_118 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_118 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3691 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3690 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3689 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3688 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3687 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3686 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3685 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3684 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3683 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3682 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3681 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3680 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3679 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3678 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3677 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3676 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3675 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3674 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3673 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3672 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3671 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3670 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3669 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3668 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3667 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3666 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3665 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3664 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3663 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3662 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3661 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV8 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV0P5SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_117 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3660 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3659 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3658 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3657 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3656 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3655 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3654 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3653 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3652 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3651 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3650 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3649 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3648 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3647 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3646 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3645 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3644 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3643 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3642 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3641 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3640 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3639 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3638 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3637 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3636 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3635 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3634 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3633 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3632 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3631 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_INHSV2SR U2 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_XOR2HSV2 U5 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_3630 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module row_other_117 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_117 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3660 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3659 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3658 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3657 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3656 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3655 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3654 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3653 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3652 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3651 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3650 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3649 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3648 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3647 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3646 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3645 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3644 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3643 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3642 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3641 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3640 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3639 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3638 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3637 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3636 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3635 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3634 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3633 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3632 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3631 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3630 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV4SR U1 ( .I(t_m_1_in), .ZN(n2) );
  LVT_CLKNHSV10 U2 ( .I(n2), .ZN(n3) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
endmodule


module cell_2_116 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3629 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3628 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3627 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3626 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3625 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3624 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3623 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3622 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3621 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3620 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3619 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3618 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3617 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3616 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3615 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3614 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3613 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3612 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3611 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3610 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3609 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3608 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3607 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3606 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3605 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3604 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3603 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3602 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV2 U5 ( .I(n6), .ZN(n4) );
  LVT_CLKXOR2HSV2 U6 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_3_3601 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3600 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3599 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_116 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4, n5;

  cell_2_116 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3629 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3628 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3627 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3626 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3625 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3624 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3623 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3622 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3621 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3620 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3619 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3618 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3617 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3616 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3615 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3614 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3613 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3612 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3611 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3610 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3609 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3608 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3607 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3606 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3605 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3604 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3603 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3602 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3601 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3600 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3599 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV1 U1 ( .I(t_m_1_in), .ZN(n3) );
  LVT_INHSV2 U2 ( .I(n3), .ZN(n4) );
  LVT_CLKNHSV5 U3 ( .I(n4), .ZN(n1) );
  LVT_INHSV10SR U4 ( .I(n1), .ZN(n2) );
  LVT_CLKNHSV4 U5 ( .I(n3), .ZN(n5) );
endmodule


module cell_2_115 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3598 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3597 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3596 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3595 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3594 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3593 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3592 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3591 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3590 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3589 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3588 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3587 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3586 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3585 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3584 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3583 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3582 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3581 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3580 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3579 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3578 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3577 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3576 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3575 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0P5 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV0SR U5 ( .I(n10), .ZN(n4) );
  LVT_CLKNHSV2 U6 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV0 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_XOR2HSV2 U8 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
endmodule


module cell_3_3574 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3573 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3572 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3571 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n5), .A2(n6), .Z(t_i_out) );
endmodule


module cell_3_3570 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3569 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3568 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_CLKNAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module row_other_115 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_115 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_3598 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3597 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3596 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3595 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3594 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3593 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3592 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3591 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3590 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3589 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3588 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3587 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3586 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3585 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3584 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3583 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3582 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3581 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3580 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3579 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3578 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3577 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3576 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3575 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3574 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3573 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3572 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3571 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3570 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3569 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3568 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_114 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_3567 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3566 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3565 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3564 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3563 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3562 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3561 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3560 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3559 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3558 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3557 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3556 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3555 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3554 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3553 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3552 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3551 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3550 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3549 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3548 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3547 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3546 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3545 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3544 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3543 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV1 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_3542 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3541 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV1 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3540 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3539 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3538 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0SR U5 ( .I(n8), .ZN(n4) );
  LVT_INHSV2 U6 ( .I(t_i_1_in), .ZN(n5) );
  LVT_CLKXOR2HSV2 U7 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV0 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_3537 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKXOR2HSV2 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module row_other_114 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_114 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3567 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3566 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3565 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3564 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3563 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3562 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3561 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3560 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3559 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3558 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3557 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3556 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3555 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3554 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3553 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3552 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3551 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3550 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3549 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3548 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3547 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3546 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3545 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3544 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3543 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3542 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3541 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3540 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3539 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3538 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3537 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV8SR U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV4 U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_113 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3536 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3535 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3534 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3533 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3532 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3531 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3530 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3529 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3528 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3527 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3526 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3525 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3524 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3523 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3522 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3521 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3520 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3519 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3518 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3517 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3516 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3515 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3514 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3513 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3512 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3511 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3510 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3509 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3508 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKXOR2HSV2 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_3507 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_3506 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_OAI21HSV2 U1 ( .A1(n6), .A2(n4), .B(n2), .ZN(t_i_out) );
  LVT_CLKNAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(t_i_1_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n6), .A2(n4), .ZN(n2) );
endmodule


module row_other_113 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_113 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3536 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3535 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3534 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3533 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3532 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3531 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3530 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3529 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3528 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3527 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3526 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3525 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3524 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3523 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3522 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3521 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3520 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3519 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3518 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3517 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3516 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3515 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3514 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3513 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3512 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3511 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3510 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3509 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3508 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3507 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3506 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV4 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_112 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3505 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3504 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3503 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3502 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3501 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3500 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3499 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3498 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3497 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3496 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3495 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3494 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3493 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3492 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3491 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3490 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3489 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3488 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3487 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3486 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3485 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3484 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3483 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3482 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3481 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U4 ( .I(n6), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_3480 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3479 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3478 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module cell_3_3477 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_XOR2HSV2 U1 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_CLKNAND2HSV1 U3 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_CLKNAND2HSV1 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U5 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_CLKNHSV0 U6 ( .I(n8), .ZN(n4) );
  LVT_INHSV2 U7 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV0 U8 ( .A1(b_in), .A2(a_in), .ZN(n8) );
endmodule


module cell_3_3476 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U2 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3475 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module row_other_112 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_112 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3505 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3504 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3503 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3502 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3501 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3500 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3499 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3498 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3497 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3496 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3495 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3494 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3493 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3492 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3491 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3490 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3489 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3488 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3487 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3486 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3485 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3484 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3483 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3482 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3481 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3480 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3479 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3478 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3477 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3476 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3475 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV5 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_111 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3474 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3473 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3472 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3471 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3470 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3469 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3468 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3467 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3466 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3465 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3464 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3463 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3462 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3461 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3460 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3459 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3458 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3457 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3456 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3455 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3454 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3453 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3452 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3451 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3450 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3449 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3448 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3447 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3446 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3445 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3444 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_111 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_111 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3474 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3473 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3472 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3471 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3470 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3469 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3468 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3467 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3466 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3465 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3464 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3463 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3462 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3461 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3460 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3459 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3458 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3457 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3456 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3455 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3454 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3453 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3452 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3451 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3450 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3449 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3448 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3447 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3446 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3445 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3444 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV6 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_110 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_3443 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3442 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3441 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3440 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3439 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3438 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3437 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3436 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3435 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3434 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3433 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3432 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3431 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3430 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3429 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3428 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3427 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3426 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3425 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3424 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3423 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3422 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3421 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3420 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3419 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3418 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3417 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3416 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3415 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3414 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module cell_3_3413 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2SR U4 ( .I(n9), .ZN(n2) );
  LVT_CLKNHSV0P5 U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV0P5 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV4 U7 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV0P5 U8 ( .A1(n9), .A2(n7), .ZN(n5) );
endmodule


module row_other_110 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4, n5;

  cell_2_110 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3443 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3442 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3441 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3440 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3439 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3438 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3437 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3436 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3435 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3434 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3433 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3432 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3431 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3430 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3429 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3428 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3427 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3426 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3425 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3424 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3423 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3422 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3421 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3420 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3419 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3418 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3417 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3416 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3415 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3414 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3413 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV2 U1 ( .I(n4), .ZN(n5) );
  LVT_INHSV2 U2 ( .I(n2), .ZN(n1) );
  LVT_INHSV0SR U3 ( .I(n5), .ZN(n2) );
  LVT_INHSV2 U4 ( .I(n2), .ZN(n3) );
  LVT_INHSV0SR U5 ( .I(t_m_1_in), .ZN(n4) );
endmodule


module cell_2_109 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_3412 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3411 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3410 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3409 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3408 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3407 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3406 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3405 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3404 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3403 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3402 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3401 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3400 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3399 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3398 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3397 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3396 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3395 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3394 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3393 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3392 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3391 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3390 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3389 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3388 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3387 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3386 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3385 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3384 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV4 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3383 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_INHSV2SR U4 ( .I(n10), .ZN(n4) );
  LVT_NAND2HSV2 U5 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U6 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_CLKNHSV2 U7 ( .I(n9), .ZN(n5) );
  LVT_CLKNAND2HSV3 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_3382 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_OAI21HSV2 U1 ( .A1(n6), .A2(n4), .B(n2), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U4 ( .A1(n6), .A2(n4), .ZN(n2) );
  LVT_XNOR2HSV4 U5 ( .A1(n5), .A2(t_i_1_in), .ZN(n4) );
endmodule


module row_other_109 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_109 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3412 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3411 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3410 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3409 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3408 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3407 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3406 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3405 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3404 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3403 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3402 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3401 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3400 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3399 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3398 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3397 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3396 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3395 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3394 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3393 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3392 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3391 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3390 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3389 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3388 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3387 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3386 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3385 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3384 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3383 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3382 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV8 U1 ( .I(n3), .ZN(n1) );
  LVT_INHSV2P5 U2 ( .I(n3), .ZN(n2) );
  LVT_CLKNHSV6 U3 ( .I(t_m_1_in), .ZN(n3) );
endmodule


module cell_2_108 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3381 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3380 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3379 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3378 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3377 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3376 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3375 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3374 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3373 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3372 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3371 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3370 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3369 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3368 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3367 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3366 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3365 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3364 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3363 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3362 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3361 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3360 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3359 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3358 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3357 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3356 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3355 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3354 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3353 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3352 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3351 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_108 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_108 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3381 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3380 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3379 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3378 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3377 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3376 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3375 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3374 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3373 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3372 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3371 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3370 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3369 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3368 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3367 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3366 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3365 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3364 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3363 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3362 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3361 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3360 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3359 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3358 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3357 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3356 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3355 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3354 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3353 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3352 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3351 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV4SR U1 ( .I(n2), .ZN(n3) );
  LVT_INHSV2 U2 ( .I(t_m_1_in), .ZN(n2) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
endmodule


module cell_2_107 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_3350 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3349 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3348 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3347 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3346 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3345 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3344 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3343 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3342 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3341 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3340 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3339 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3338 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3337 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3336 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3335 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3334 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3333 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3332 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3331 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3330 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3329 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3328 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3327 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3326 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3325 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3324 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3323 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3322 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3321 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_CLKNAND2HSV1 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV0 U4 ( .I(n6), .ZN(n4) );
  LVT_XOR2HSV2 U5 ( .A1(n7), .A2(n8), .Z(t_i_out) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_3320 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV4 U2 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_CLKAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .Z(n3) );
  LVT_XNOR2HSV4 U4 ( .A1(n3), .A2(t_i_1_in), .ZN(n4) );
endmodule


module row_other_107 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_2_107 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3350 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3349 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3348 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3347 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3346 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3345 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3344 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3343 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3342 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3341 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3340 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3339 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3338 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3337 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3336 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3335 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3334 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3333 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3332 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3331 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3330 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3329 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3328 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3327 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3326 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3325 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3324 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3323 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3322 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3321 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3320 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV4SR U1 ( .I(n3), .ZN(n4) );
  LVT_INHSV2SR U2 ( .I(t_m_1_in), .ZN(n3) );
  LVT_INHSV0SR U3 ( .I(n4), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_106 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3319 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3318 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3317 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3316 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3315 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3314 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3313 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3312 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3311 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3310 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3309 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3308 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3307 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3306 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3305 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3304 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3303 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3302 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3301 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3300 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3299 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3298 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3297 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3296 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3295 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3294 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3293 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3292 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3291 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_CLKXOR2HSV2 U1 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV4 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U3 ( .A1(n3), .A2(t_i_1_in), .ZN(n4) );
  LVT_CLKAND2HSV2 U4 ( .A1(b_in), .A2(a_in), .Z(n3) );
endmodule


module cell_3_3290 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_3289 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_106 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_106 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3319 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3318 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3317 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3316 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3315 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3314 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3313 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3312 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3311 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3310 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3309 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3308 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3307 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3306 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3305 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3304 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3303 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3302 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3301 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3300 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3299 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3298 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3297 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3296 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3295 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3294 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3293 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3292 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3291 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3290 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3289 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV6 U1 ( .I(n2), .ZN(n3) );
  LVT_INHSV2 U2 ( .I(t_m_1_in), .ZN(n2) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
endmodule


module cell_2_105 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3288 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3287 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3286 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3285 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3284 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3283 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3282 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3281 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3280 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3279 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3278 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3277 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3276 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3275 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3274 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3273 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3272 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3271 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3270 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3269 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3268 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3267 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3266 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3265 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3264 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3263 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_XOR2HSV0 U1 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV0P5 U2 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0 U3 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U5 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0SR U6 ( .I(n8), .ZN(n4) );
  LVT_CLKNHSV2 U7 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV2 U8 ( .A1(b_in), .A2(a_in), .ZN(n8) );
endmodule


module cell_3_3262 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3261 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3260 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3259 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_INHSV2 U2 ( .I(n8), .ZN(n4) );
  LVT_XOR2HSV4 U4 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_OAI21HSV2 U6 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
endmodule


module cell_3_3258 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV8 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_105 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_105 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_3288 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3287 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3286 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3285 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3284 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3283 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3282 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3281 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3280 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3279 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3278 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3277 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3276 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3275 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3274 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3273 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3272 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3271 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3270 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3269 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3268 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3267 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3266 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3265 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3264 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3263 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3262 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3261 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3260 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3259 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3258 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_104 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3257 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3256 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3255 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3254 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3253 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3252 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3251 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3250 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3249 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3248 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3247 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3246 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3245 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3244 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3243 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3242 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3241 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3240 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3239 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3238 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3237 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3236 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3235 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3234 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3233 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3232 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3231 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3230 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV2 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_3229 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3228 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3227 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module row_other_104 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_104 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3257 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3256 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3255 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3254 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3253 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3252 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3251 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3250 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3249 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3248 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3247 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3246 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3245 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3244 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3243 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3242 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3241 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3240 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3239 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3238 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3237 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3236 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3235 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3234 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3233 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3232 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3231 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3230 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3229 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3228 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3227 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2 U1 ( .I(t_m_1_in), .ZN(n2) );
  LVT_INHSV4 U2 ( .I(n2), .ZN(n1) );
endmodule


module cell_2_103 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_3226 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3225 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3224 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3223 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3222 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3221 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3220 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3219 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3218 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3217 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3216 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3215 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3214 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3213 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3212 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3211 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3210 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3209 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3208 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3207 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3206 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3205 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3204 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3203 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3202 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3201 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3200 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3199 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_3198 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_NAND2HSV0P5 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_CLKXOR2HSV4 U2 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U5 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV2 U6 ( .I(n8), .ZN(n4) );
  LVT_INHSV2 U7 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV0 U8 ( .A1(b_in), .A2(a_in), .ZN(n8) );
endmodule


module cell_3_3197 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3196 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNHSV2 U1 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV1 U2 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV4 U5 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U8 ( .I(n7), .ZN(n4) );
endmodule


module row_other_103 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_103 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3226 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3225 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3224 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3223 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3222 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3221 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3220 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3219 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3218 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3217 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3216 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3215 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3214 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3213 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3212 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3211 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3210 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3209 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3208 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3207 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3206 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3205 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3204 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3203 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3202 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3201 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3200 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3199 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3198 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3197 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3196 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV1SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_CLKNHSV4 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_102 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3195 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3194 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3193 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3192 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3191 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3190 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3189 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3188 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3187 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3186 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3185 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3184 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3183 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3182 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3181 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3180 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3179 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3178 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3177 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3176 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3175 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3174 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3173 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3172 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3171 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3170 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3169 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3168 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3167 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n9), .A2(n5), .ZN(n6) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n4), .A2(n10), .ZN(n7) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV2SR U5 ( .I(n9), .ZN(n4) );
  LVT_INHSV2P5 U6 ( .I(n10), .ZN(n5) );
  LVT_XOR2HSV2 U7 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_NAND2HSV0P5 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_3166 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_CLKNHSV2 U1 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV2 U3 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV2 U5 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U6 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U7 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV2 U8 ( .I(n8), .ZN(n4) );
endmodule


module cell_3_3165 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV2 U1 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_INHSV2 U5 ( .I(n7), .ZN(n4) );
  LVT_INHSV1SR U6 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV0P5 U7 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_102 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_102 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3195 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3194 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3193 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3192 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3191 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3190 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3189 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3188 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3187 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3186 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3185 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3184 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3183 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3182 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3181 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3180 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3179 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3178 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3177 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3176 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3175 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3174 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3173 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3172 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3171 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3170 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3169 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3168 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3167 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3166 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3165 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2 U1 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U2 ( .I(t_m_1_in), .ZN(n3) );
  LVT_INHSV4SR U3 ( .I(n3), .ZN(n1) );
endmodule


module cell_2_101 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_3164 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3163 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3162 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3161 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3160 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3159 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3158 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3157 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3156 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3155 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3154 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3153 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3152 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3151 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3150 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3149 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3148 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3147 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3146 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3145 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3144 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3143 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3142 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3141 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3140 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3139 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV3 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3138 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3137 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3136 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3135 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_3134 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV1 U1 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV0P5SR U2 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV4 U5 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV4 U6 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV4 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_101 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_101 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3164 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3163 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3162 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3161 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3160 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3159 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3158 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3157 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3156 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3155 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3154 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3153 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3152 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3151 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3150 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3149 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3148 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3147 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3146 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3145 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3144 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3143 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3142 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3141 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3140 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3139 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3138 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3137 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3136 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3135 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3134 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2SR U1 ( .I(t_m_1_in), .ZN(n2) );
  LVT_CLKNHSV4 U2 ( .I(n2), .ZN(n1) );
endmodule


module cell_2_100 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_3133 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3132 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3131 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3130 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3129 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3128 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3127 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3126 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3125 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3124 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3123 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3122 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3121 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3120 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3119 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3118 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3117 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3116 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3115 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3114 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3113 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3112 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3111 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3110 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3109 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U3 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U5 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_3_3108 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3107 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3106 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(n5), .A2(n6), .Z(t_i_out) );
endmodule


module cell_3_3105 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3104 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3103 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_100 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1;

  cell_2_100 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_3133 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3132 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3131 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3130 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3129 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3128 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3127 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3126 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3125 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3124 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3123 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3122 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3121 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3120 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3119 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3118 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3117 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3116 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3115 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3114 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3113 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3112 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3111 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3110 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3109 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3108 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3107 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3106 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3105 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3104 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3103 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV4 U1 ( .I(t_m_1_in), .Z(n1) );
endmodule


module cell_2_99 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3102 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3101 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3100 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3099 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3098 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3097 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3096 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3095 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3094 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3093 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3092 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3091 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3090 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3089 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3088 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3087 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3086 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3085 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3084 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3083 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3082 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3081 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3080 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3079 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3078 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3077 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3076 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3075 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3074 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3073 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3072 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n9) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n2), .A2(n4), .ZN(n5) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n5), .A2(n7), .ZN(t_i_out) );
  LVT_CLKNHSV2 U4 ( .I(n6), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV4 U6 ( .A1(n10), .A2(n8), .ZN(n7) );
  LVT_NAND2HSV0 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(n9), .A2(t_i_1_in), .ZN(n8) );
  LVT_NAND2HSV2 U9 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module row_other_99 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_99 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_3102 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3101 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3100 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3099 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3098 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3097 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3096 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3095 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3094 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3093 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3092 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3091 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3090 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3089 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3088 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3087 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3086 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3085 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3084 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3083 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3082 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3081 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3080 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3079 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3078 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3077 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3076 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3075 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3074 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3073 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3072 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_98 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3071 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3070 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3069 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3068 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3067 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3066 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3065 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3064 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3063 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3062 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3061 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3060 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3059 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3058 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3057 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3056 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3055 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3054 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3053 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3052 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3051 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3050 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3049 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3048 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3047 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3046 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3045 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3044 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3043 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3042 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3041 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_98 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_98 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_3071 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3070 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3069 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3068 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3067 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3066 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3065 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3064 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3063 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3062 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3061 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3060 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3059 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3058 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3057 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3056 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3055 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3054 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3053 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3052 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3051 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3050 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3049 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3048 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3047 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3046 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3045 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3044 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3043 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3042 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3041 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV4 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV2SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_97 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_3040 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3039 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3038 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3037 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3036 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3035 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3034 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3033 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3032 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3031 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3030 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3029 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3028 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3027 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3026 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3025 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3024 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3023 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3022 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3021 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3020 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3019 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3018 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3017 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3016 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3015 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3014 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3013 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3012 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3011 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3010 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_CLKNAND2HSV1 U1 ( .A1(n6), .A2(n8), .ZN(n4) );
  LVT_NAND2HSV8 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n5), .A2(n4), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U5 ( .A1(n7), .A2(t_i_1_in), .ZN(n6) );
  LVT_INAND2HSV4 U6 ( .A1(n8), .B1(n2), .ZN(n5) );
  LVT_INHSV2 U7 ( .I(n6), .ZN(n2) );
endmodule


module row_other_97 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_2_97 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_3040 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3039 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3038 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3037 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3036 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3035 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3034 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3033 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3032 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3031 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_3030 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_3029 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_3028 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_3027 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_3026 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_3025 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_3024 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_3023 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_3022 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_3021 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_3020 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_3019 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_3018 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_3017 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_3016 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_3015 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_3014 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3013 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_3012 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_3011 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_3010 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV12SR U1 ( .I(n1), .ZN(n3) );
  LVT_INHSV2P5 U2 ( .I(n1), .ZN(n4) );
  LVT_INHSV6 U3 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2SR U4 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_96 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_3009 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_3008 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3007 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3006 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3005 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3004 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3003 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3002 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3001 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_3000 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2999 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2998 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2997 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2996 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2995 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2994 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2993 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2992 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2991 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2990 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2989 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2988 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2987 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2986 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2985 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2984 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2983 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2982 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_2981 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2980 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_2979 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U4 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV4 U5 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2 U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV1 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_96 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_96 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_3009 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_3008 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_3007 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_3006 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_3005 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_3004 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_3003 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_3002 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_3001 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_3000 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2999 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2998 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2997 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2996 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2995 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2994 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2993 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2992 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2991 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2990 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2989 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2988 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2987 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2986 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2985 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2984 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2983 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2982 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2981 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2980 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2979 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_95 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_2978 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2977 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2976 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2975 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2974 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2973 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2972 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2971 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2970 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2969 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2968 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2967 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2966 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2965 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2964 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2963 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2962 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2961 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2960 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2959 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2958 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2957 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2956 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2955 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2954 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2953 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2952 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2951 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2950 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2949 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2948 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_OAI21HSV2 U1 ( .A1(t_i_1_in), .A2(n5), .B(n2), .ZN(n4) );
  LVT_CLKNAND2HSV1 U2 ( .A1(n5), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV12 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_NAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_XNOR2HSV4 U5 ( .A1(n6), .A2(n4), .ZN(t_i_out) );
endmodule


module row_other_95 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_95 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_2978 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2977 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2976 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2975 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2974 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2973 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2972 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2971 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2970 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2969 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2968 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2967 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2966 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2965 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2964 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2963 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2962 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2961 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2960 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2959 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2958 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2957 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2956 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2955 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2954 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2953 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2952 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2951 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2950 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2949 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2948 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_94 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_2947 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2946 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2945 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2944 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2943 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2942 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2941 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2940 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2939 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2938 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2937 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2936 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2935 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2934 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2933 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2932 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2931 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2930 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2929 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2928 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2927 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2926 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2925 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2924 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2923 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2922 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2921 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2920 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2919 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2918 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2917 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV4 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV2 U2 ( .I(n7), .ZN(n4) );
  LVT_CLKNHSV2 U4 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV2 U5 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV4 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_94 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_94 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_2947 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2946 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2945 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2944 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2943 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2942 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2941 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2940 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2939 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2938 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2937 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2936 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2935 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2934 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2933 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2932 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2931 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2930 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2929 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2928 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2927 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2926 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2925 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2924 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2923 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2922 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2921 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2920 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2919 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2918 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2917 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_93 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4, n5, n6;

  LVT_OAI21HSV1 U1 ( .A1(n3), .A2(n5), .B(n4), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_NAND2HSV0P5 U3 ( .A1(n3), .A2(n5), .ZN(n4) );
  LVT_INHSV0SR U4 ( .I(n6), .ZN(n3) );
  LVT_CLKNAND2HSV1 U5 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_3_2916 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2915 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2914 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2913 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2912 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2911 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2910 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2909 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2908 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2907 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2906 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2905 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2904 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2903 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2902 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2901 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2900 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2899 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2898 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2897 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2896 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2895 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2894 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2893 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2892 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2891 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2890 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2889 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2888 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2887 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2886 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module row_other_93 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_93 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_2916 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2915 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2914 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2913 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2912 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2911 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2910 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2909 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2908 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2907 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2906 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2905 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2904 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2903 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2902 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2901 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2900 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2899 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2898 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2897 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2896 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2895 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2894 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2893 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2892 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2891 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2890 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2889 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2888 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2887 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2886 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_3 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [31:0] a_in;
  input [31:0] g_in;
  input [31:0] b_in;
  input [31:0] t_m_1_in;
  input [30:0] t_i_1_in;
  input [30:0] t_i_2_in;
  output [31:0] a_out;
  output [31:0] g_out;
  output [30:0] t_i_1_out;
  output [30:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;
  wire   n1, n2, n4, n5, n7, n8, n10, n11, n13, n15, n16, n18, n20, n21, n23,
         n25;
  wire   [30:0] t0;
  wire   [30:0] t1;
  wire   [30:0] t2;
  wire   [30:0] t3;
  wire   [30:0] t4;
  wire   [30:0] t5;
  wire   [30:0] t6;
  wire   [30:0] t7;
  wire   [30:0] t8;
  wire   [30:0] t9;
  wire   [30:0] t10;
  wire   [30:0] t11;
  wire   [30:0] t12;
  wire   [30:0] t13;
  wire   [30:0] t14;
  wire   [30:0] t15;
  wire   [30:0] t16;
  wire   [30:0] t17;
  wire   [30:0] t18;
  wire   [30:0] t19;
  wire   [30:0] t20;
  wire   [30:0] t21;
  wire   [30:0] t22;
  wire   [30:0] t23;
  wire   [30:0] t24;
  wire   [30:0] t25;
  wire   [30:0] t26;
  wire   [30:0] t27;
  wire   [30:0] t28;
  wire   [30:0] t29;
  wire   [30:0] t30;
  assign a_out[31] = a_in[31];
  assign a_out[29] = a_in[29];
  assign a_out[23] = a_in[23];
  assign a_out[22] = a_in[22];
  assign a_out[21] = a_in[21];
  assign a_out[20] = a_in[20];
  assign a_out[19] = a_in[19];
  assign a_out[18] = a_in[18];
  assign a_out[17] = a_in[17];
  assign a_out[16] = a_in[16];
  assign a_out[15] = a_in[15];
  assign a_out[14] = a_in[14];
  assign a_out[13] = a_in[13];
  assign a_out[12] = a_in[12];
  assign a_out[11] = a_in[11];
  assign a_out[10] = a_in[10];
  assign a_out[9] = a_in[9];
  assign a_out[8] = a_in[8];
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[31] = g_in[31];
  assign g_out[30] = g_in[30];
  assign g_out[28] = g_in[28];
  assign g_out[27] = g_in[27];
  assign g_out[23] = g_in[23];
  assign g_out[22] = g_in[22];
  assign g_out[21] = g_in[21];
  assign g_out[20] = g_in[20];
  assign g_out[19] = g_in[19];
  assign g_out[18] = g_in[18];
  assign g_out[17] = g_in[17];
  assign g_out[16] = g_in[16];
  assign g_out[15] = g_in[15];
  assign g_out[14] = g_in[14];
  assign g_out[13] = g_in[13];
  assign g_out[12] = g_in[12];
  assign g_out[11] = g_in[11];
  assign g_out[10] = g_in[10];
  assign g_out[9] = g_in[9];
  assign g_out[8] = g_in[8];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_3 u0 ( .a_in({a_in[31:28], n21, n16, n5, a_in[24:0]}), .g_in({
        g_in[31:30], n8, g_in[28:27], n13, n2, n11, g_in[23:0]}), .b_in(
        b_in[31]), .t_m_1_in(t_m_1_in[31]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), 
        .t_i_2_in(t_i_2_in), .t_i_1_out(t0), .t_i_2_out(t_i_2_out[30]) );
  row_other_123 u1 ( .a_in({a_in[31:29], a_out[28:24], a_in[23:0]}), .g_in({
        g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], g_in[23:0]}), 
        .b_in(b_in[30]), .t_m_1_in(t_m_1_in[30]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(t_i_2_out[29]) );
  row_other_122 u2 ( .a_in({a_in[31:29], a_out[28:24], a_in[23:0]}), .g_in({
        g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], g_in[23:0]}), 
        .b_in(b_in[29]), .t_m_1_in(t_m_1_in[29]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(t_i_2_out[28]) );
  row_other_121 u3 ( .a_in({a_in[31:29], a_out[28:24], a_in[23:0]}), .g_in({
        g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], g_in[23:0]}), 
        .b_in(b_in[28]), .t_m_1_in(t_m_1_in[28]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(t_i_2_out[27]) );
  row_other_120 u4 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[27]), .t_m_1_in(t_m_1_in[27]), .t_i_1_in(t3), 
        .t_i_1_out(t4), .t_i_2_out(t_i_2_out[26]) );
  row_other_119 u5 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[26]), .t_m_1_in(t_m_1_in[26]), .t_i_1_in(t4), 
        .t_i_1_out(t5), .t_i_2_out(t_i_2_out[25]) );
  row_other_118 u6 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[25]), .t_m_1_in(t_m_1_in[25]), .t_i_1_in(t5), 
        .t_i_1_out(t6), .t_i_2_out(t_i_2_out[24]) );
  row_other_117 u7 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[24]), .t_m_1_in(t_m_1_in[24]), .t_i_1_in(t6), 
        .t_i_1_out(t7), .t_i_2_out(t_i_2_out[23]) );
  row_other_116 u8 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[23]), .t_m_1_in(t_m_1_in[23]), .t_i_1_in(t7), 
        .t_i_1_out(t8), .t_i_2_out(t_i_2_out[22]) );
  row_other_115 u9 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[22]), .t_m_1_in(t_m_1_in[22]), .t_i_1_in(t8), 
        .t_i_1_out(t9), .t_i_2_out(t_i_2_out[21]) );
  row_other_114 u10 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[21]), .t_m_1_in(t_m_1_in[21]), .t_i_1_in(t9), 
        .t_i_1_out(t10), .t_i_2_out(t_i_2_out[20]) );
  row_other_113 u11 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[20]), .t_m_1_in(t_m_1_in[20]), .t_i_1_in(t10), 
        .t_i_1_out(t11), .t_i_2_out(t_i_2_out[19]) );
  row_other_112 u12 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[19]), .t_m_1_in(t_m_1_in[19]), .t_i_1_in(t11), 
        .t_i_1_out(t12), .t_i_2_out(t_i_2_out[18]) );
  row_other_111 u13 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[18]), .t_m_1_in(t_m_1_in[18]), .t_i_1_in(t12), 
        .t_i_1_out(t13), .t_i_2_out(t_i_2_out[17]) );
  row_other_110 u14 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[17]), .t_m_1_in(t_m_1_in[17]), .t_i_1_in(t13), 
        .t_i_1_out(t14), .t_i_2_out(t_i_2_out[16]) );
  row_other_109 u15 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[16]), .t_m_1_in(t_m_1_in[16]), .t_i_1_in(t14), 
        .t_i_1_out(t15), .t_i_2_out(t_i_2_out[15]) );
  row_other_108 u16 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[15]), .t_m_1_in(t_m_1_in[15]), .t_i_1_in(t15), 
        .t_i_1_out(t16), .t_i_2_out(t_i_2_out[14]) );
  row_other_107 u17 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[14]), .t_m_1_in(t_m_1_in[14]), .t_i_1_in(t16), 
        .t_i_1_out(t17), .t_i_2_out(t_i_2_out[13]) );
  row_other_106 u18 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[13]), .t_m_1_in(t_m_1_in[13]), .t_i_1_in(t17), 
        .t_i_1_out(t18), .t_i_2_out(t_i_2_out[12]) );
  row_other_105 u19 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[12]), .t_m_1_in(t_m_1_in[12]), .t_i_1_in(t18), 
        .t_i_1_out(t19), .t_i_2_out(t_i_2_out[11]) );
  row_other_104 u20 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[11]), .t_m_1_in(t_m_1_in[11]), .t_i_1_in(t19), 
        .t_i_1_out(t20), .t_i_2_out(t_i_2_out[10]) );
  row_other_103 u21 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[10]), .t_m_1_in(t_m_1_in[10]), .t_i_1_in(t20), 
        .t_i_1_out(t21), .t_i_2_out(t_i_2_out[9]) );
  row_other_102 u22 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[9]), .t_m_1_in(t_m_1_in[9]), .t_i_1_in(t21), 
        .t_i_1_out(t22), .t_i_2_out(t_i_2_out[8]) );
  row_other_101 u23 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[8]), .t_m_1_in(t_m_1_in[8]), .t_i_1_in(t22), 
        .t_i_1_out(t23), .t_i_2_out(t_i_2_out[7]) );
  row_other_100 u24 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[7]), .t_m_1_in(t_m_1_in[7]), .t_i_1_in(t23), 
        .t_i_1_out(t24), .t_i_2_out(t_i_2_out[6]) );
  row_other_99 u25 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[6]), .t_m_1_in(t_m_1_in[6]), .t_i_1_in(t24), 
        .t_i_1_out(t25), .t_i_2_out(t_i_2_out[5]) );
  row_other_98 u26 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[5]), .t_m_1_in(t_m_1_in[5]), .t_i_1_in(t25), 
        .t_i_1_out(t26), .t_i_2_out(t_i_2_out[4]) );
  row_other_97 u27 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[4]), .t_m_1_in(t_m_1_in[4]), .t_i_1_in(t26), 
        .t_i_1_out(t27), .t_i_2_out(t_i_2_out[3]) );
  row_other_96 u28 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[3]), .t_m_1_in(t_m_1_in[3]), .t_i_1_in(t27), 
        .t_i_1_out(t28), .t_i_2_out(t_i_2_out[2]) );
  row_other_95 u29 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[2]), .t_m_1_in(t_m_1_in[2]), .t_i_1_in(t28), 
        .t_i_1_out(t29), .t_i_2_out(t_i_2_out[1]) );
  row_other_94 u30 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[1]), .t_m_1_in(t_m_1_in[1]), .t_i_1_in(t29), 
        .t_i_1_out(t30), .t_i_2_out(t_i_2_out[0]) );
  row_other_93 u31 ( .a_in({a_in[31], a_out[30], a_in[29], a_out[28:24], 
        a_in[23:0]}), .g_in({g_in[31:30], g_out[29], g_in[28:27], g_out[26:24], 
        g_in[23:0]}), .b_in(b_in[0]), .t_m_1_in(t_m_1_in[0]), .t_i_1_in(t30), 
        .t_i_1_out(t_i_1_out), .t_i_2_out(t_i_1_out_0) );
  LVT_CLKNHSV4 U1 ( .I(g_in[25]), .ZN(n1) );
  LVT_INHSV2SR U2 ( .I(n1), .ZN(n2) );
  LVT_INHSV2SR U3 ( .I(n1), .ZN(g_out[25]) );
  LVT_CLKNHSV4 U4 ( .I(a_in[25]), .ZN(n4) );
  LVT_INHSV2SR U5 ( .I(n4), .ZN(n5) );
  LVT_INHSV2SR U6 ( .I(n4), .ZN(a_out[25]) );
  LVT_CLKNHSV2P5 U7 ( .I(g_in[29]), .ZN(n7) );
  LVT_INHSV2SR U8 ( .I(n7), .ZN(n8) );
  LVT_INHSV2SR U9 ( .I(n7), .ZN(g_out[29]) );
  LVT_CLKNHSV5 U10 ( .I(g_in[24]), .ZN(n10) );
  LVT_INHSV3SR U11 ( .I(n10), .ZN(n11) );
  LVT_INHSV2SR U12 ( .I(n10), .ZN(g_out[24]) );
  LVT_BUFHSV2 U13 ( .I(g_in[26]), .Z(n13) );
  LVT_INHSV2 U14 ( .I(a_in[26]), .ZN(n15) );
  LVT_BUFHSV2RT U15 ( .I(g_in[26]), .Z(g_out[26]) );
  LVT_INHSV2SR U16 ( .I(n15), .ZN(n16) );
  LVT_INHSV2SR U17 ( .I(n15), .ZN(a_out[26]) );
  LVT_INHSV2 U18 ( .I(a_in[27]), .ZN(n20) );
  LVT_INHSV2 U19 ( .I(a_in[24]), .ZN(n18) );
  LVT_INHSV2 U20 ( .I(a_in[28]), .ZN(n23) );
  LVT_INHSV2SR U21 ( .I(n18), .ZN(a_out[24]) );
  LVT_INHSV2SR U22 ( .I(n20), .ZN(n21) );
  LVT_INHSV2SR U23 ( .I(n20), .ZN(a_out[27]) );
  LVT_INHSV2SR U24 ( .I(n23), .ZN(a_out[28]) );
  LVT_INHSV0SR U25 ( .I(a_in[30]), .ZN(n25) );
  LVT_INHSV2 U26 ( .I(n25), .ZN(a_out[30]) );
endmodule


module regist_32bit_19 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_32bit_18 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_31bit_12 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module PE_3 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro );
  input [31:0] a_in;
  input [31:0] g_in;
  input [31:0] b_in;
  input [30:0] t_i_1_in;
  input [30:0] t_i_2_in;
  output [31:0] a_out;
  output [31:0] g_out;
  output [31:0] b_out;
  output [30:0] t_i_1_out;
  output [30:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0, to_1, ti_1, n2,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94;
  wire   [31:0] l_a;
  wire   [31:0] l_g;
  wire   [30:0] l_t_i_1_in;
  wire   [30:0] l_t_i_2_in;
  wire   [31:0] mux_b;
  wire   [31:0] mux_bq;
  wire   [30:0] to_7;
  wire   [30:0] ti_7;
  wire   [31:0] ao;
  wire   [31:0] go;
  wire   [30:0] to;

  LVT_AO22HSV0 U35 ( .A1(mux_bq[9]), .A2(n58), .B1(b_out[9]), .B2(n34), .Z(
        mux_b[9]) );
  LVT_AO22HSV0 U36 ( .A1(mux_bq[8]), .A2(n58), .B1(b_out[8]), .B2(n34), .Z(
        mux_b[8]) );
  LVT_AO22HSV0 U37 ( .A1(mux_bq[7]), .A2(n58), .B1(b_out[7]), .B2(n34), .Z(
        mux_b[7]) );
  LVT_AO22HSV0 U38 ( .A1(mux_bq[6]), .A2(n58), .B1(b_out[6]), .B2(n34), .Z(
        mux_b[6]) );
  LVT_AO22HSV0 U39 ( .A1(mux_bq[5]), .A2(n58), .B1(b_out[5]), .B2(n34), .Z(
        mux_b[5]) );
  LVT_AO22HSV0 U40 ( .A1(mux_bq[4]), .A2(n58), .B1(b_out[4]), .B2(n34), .Z(
        mux_b[4]) );
  LVT_AO22HSV0 U41 ( .A1(mux_bq[3]), .A2(n58), .B1(b_out[3]), .B2(n34), .Z(
        mux_b[3]) );
  LVT_AO22HSV0 U42 ( .A1(n30), .A2(n58), .B1(b_out[31]), .B2(n34), .Z(
        mux_b[31]) );
  LVT_AO22HSV0 U43 ( .A1(mux_bq[30]), .A2(n58), .B1(b_out[30]), .B2(n34), .Z(
        mux_b[30]) );
  LVT_AO22HSV0 U44 ( .A1(mux_bq[2]), .A2(n58), .B1(b_out[2]), .B2(n34), .Z(
        mux_b[2]) );
  LVT_AO22HSV0 U45 ( .A1(mux_bq[29]), .A2(n58), .B1(b_out[29]), .B2(n34), .Z(
        mux_b[29]) );
  LVT_AO22HSV0 U46 ( .A1(mux_bq[28]), .A2(n58), .B1(b_out[28]), .B2(n34), .Z(
        mux_b[28]) );
  LVT_AO22HSV0 U47 ( .A1(mux_bq[27]), .A2(n58), .B1(b_out[27]), .B2(n34), .Z(
        mux_b[27]) );
  LVT_AO22HSV0 U48 ( .A1(mux_bq[26]), .A2(n58), .B1(b_out[26]), .B2(n93), .Z(
        mux_b[26]) );
  LVT_AO22HSV0 U49 ( .A1(mux_bq[25]), .A2(n58), .B1(b_out[25]), .B2(n93), .Z(
        mux_b[25]) );
  LVT_AO22HSV0 U50 ( .A1(mux_bq[24]), .A2(n58), .B1(b_out[24]), .B2(n93), .Z(
        mux_b[24]) );
  LVT_AO22HSV0 U51 ( .A1(mux_bq[23]), .A2(n58), .B1(b_out[23]), .B2(n93), .Z(
        mux_b[23]) );
  LVT_AO22HSV0 U52 ( .A1(mux_bq[22]), .A2(n58), .B1(b_out[22]), .B2(n93), .Z(
        mux_b[22]) );
  LVT_AO22HSV0 U53 ( .A1(mux_bq[21]), .A2(n58), .B1(b_out[21]), .B2(n93), .Z(
        mux_b[21]) );
  LVT_AO22HSV0 U54 ( .A1(mux_bq[20]), .A2(n58), .B1(b_out[20]), .B2(n93), .Z(
        mux_b[20]) );
  LVT_AO22HSV0 U55 ( .A1(mux_bq[1]), .A2(n58), .B1(b_out[1]), .B2(n34), .Z(
        mux_b[1]) );
  LVT_AO22HSV0 U56 ( .A1(mux_bq[19]), .A2(n58), .B1(b_out[19]), .B2(n93), .Z(
        mux_b[19]) );
  LVT_AO22HSV0 U57 ( .A1(mux_bq[18]), .A2(n58), .B1(b_out[18]), .B2(n93), .Z(
        mux_b[18]) );
  LVT_AO22HSV0 U58 ( .A1(mux_bq[17]), .A2(n58), .B1(b_out[17]), .B2(n93), .Z(
        mux_b[17]) );
  LVT_AO22HSV0 U59 ( .A1(mux_bq[16]), .A2(n58), .B1(b_out[16]), .B2(n93), .Z(
        mux_b[16]) );
  LVT_AO22HSV0 U60 ( .A1(mux_bq[15]), .A2(n58), .B1(b_out[15]), .B2(n93), .Z(
        mux_b[15]) );
  LVT_AO22HSV0 U61 ( .A1(mux_bq[14]), .A2(n58), .B1(b_out[14]), .B2(n93), .Z(
        mux_b[14]) );
  LVT_AO22HSV0 U62 ( .A1(mux_bq[13]), .A2(n58), .B1(b_out[13]), .B2(n93), .Z(
        mux_b[13]) );
  LVT_AO22HSV0 U63 ( .A1(mux_bq[12]), .A2(n58), .B1(b_out[12]), .B2(n93), .Z(
        mux_b[12]) );
  LVT_AO22HSV0 U64 ( .A1(mux_bq[11]), .A2(n58), .B1(b_out[11]), .B2(n34), .Z(
        mux_b[11]) );
  LVT_AO22HSV0 U65 ( .A1(mux_bq[10]), .A2(n58), .B1(b_out[10]), .B2(n34), .Z(
        mux_b[10]) );
  LVT_AO22HSV0 U66 ( .A1(mux_bq[0]), .A2(n58), .B1(b_out[0]), .B2(n34), .Z(
        mux_b[0]) );
  LVT_AOI21HSV0 U69 ( .A1(n92), .A2(n91), .B(n93), .ZN(\c_t_i_1_in[0] ) );
  LVT_AND4HSV0 U71 ( .A1(n90), .A2(n89), .A3(n88), .A4(n87), .Z(n91) );
  LVT_NOR4HSV0 U72 ( .A1(l_t_i_1_in[9]), .A2(l_t_i_1_in[8]), .A3(l_t_i_1_in[7]), .A4(l_t_i_1_in[6]), .ZN(n87) );
  LVT_NOR4HSV0 U73 ( .A1(l_t_i_1_in[5]), .A2(l_t_i_1_in[4]), .A3(l_t_i_1_in[3]), .A4(l_t_i_1_in[30]), .ZN(n88) );
  LVT_NOR4HSV0 U74 ( .A1(l_t_i_1_in[2]), .A2(l_t_i_1_in[29]), .A3(
        l_t_i_1_in[28]), .A4(l_t_i_1_in[27]), .ZN(n89) );
  LVT_NOR4HSV0 U75 ( .A1(l_t_i_1_in[26]), .A2(l_t_i_1_in[25]), .A3(
        l_t_i_1_in[24]), .A4(l_t_i_1_in[23]), .ZN(n90) );
  LVT_AND4HSV0 U76 ( .A1(n86), .A2(n85), .A3(n84), .A4(n83), .Z(n92) );
  LVT_NOR4HSV0 U77 ( .A1(l_t_i_1_in[22]), .A2(l_t_i_1_in[21]), .A3(
        l_t_i_1_in[20]), .A4(l_t_i_1_in[1]), .ZN(n83) );
  LVT_NOR4HSV0 U78 ( .A1(l_t_i_1_in[19]), .A2(l_t_i_1_in[18]), .A3(
        l_t_i_1_in[17]), .A4(l_t_i_1_in[16]), .ZN(n84) );
  LVT_NOR4HSV0 U79 ( .A1(l_t_i_1_in[15]), .A2(l_t_i_1_in[14]), .A3(
        l_t_i_1_in[13]), .A4(l_t_i_1_in[12]), .ZN(n85) );
  LVT_NOR3HSV0 U80 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[11]), .A3(
        l_t_i_1_in[10]), .ZN(n86) );
  regist_32bit_23 u0 ( .clk(clk), .rstn(rstn), .in(a_in), .out(l_a) );
  regist_32bit_22 u1 ( .clk(clk), .rstn(rstn), .in(b_in), .out(b_out) );
  regist_32bit_21 u2 ( .clk(clk), .rstn(rstn), .in(g_in), .out(l_g) );
  regist_1bit_15 u3 ( .clk(clk), .rstn(rstn), .in(ctr), .out(l_ctr) );
  regist_1bit_14 u4 ( .clk(clk), .rstn(rstn), .in(n58), .out(ctro) );
  regist_31bit_15 u5 ( .clk(clk), .rstn(rstn), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_31bit_14 u6 ( .clk(clk), .rstn(rstn), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_13 u7 ( .clk(clk), .rstn(rstn), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_32bit_20 u9 ( .clk(clk), .rstn(rstn), .in(mux_b), .out(mux_bq) );
  regist_1bit_12 u10 ( .clk(clk), .rstn(rstn), .in(to_1), .out(ti_1) );
  regist_31bit_13 u11 ( .clk(clk), .rstn(rstn), .in({n77, to_7[29:28], n72, 
        n66, to_7[25:21], n78, n73, n74, to_7[17:16], n33, to_7[14:13], n14, 
        to_7[11], n79, n70, to_7[8:7], n32, n75, to_7[4], n76, n18, to_7[1], 
        n67}), .out(ti_7) );
  PE_core_3 pe ( .a_in(l_a), .g_in({l_g[31:28], n22, l_g[26:25], n20, 
        l_g[23:0]}), .b_in({n30, mux_bq[30:0]}), .t_m_1_in({to_1, n77, 
        to_7[29:28], n72, n66, to_7[25:21], n78, n73, n74, to_7[17:16], n33, 
        to_7[14:11], n79, n70, to_7[8:7], n32, n75, to_7[4], n76, to_7[2:1], 
        n67}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(go), 
        .t_i_1_out(to), .t_i_2_out(t_i_2_out), .t_i_1_out_0(t_i_1_out_0) );
  regist_32bit_19 u12 ( .clk(clk), .rstn(rstn), .in(ao), .out(a_out) );
  regist_32bit_18 u13 ( .clk(clk), .rstn(rstn), .in(go), .out(g_out) );
  regist_31bit_12 u14 ( .clk(clk), .rstn(rstn), .in(to), .out(t_i_1_out) );
  LVT_CLKNAND2HSV4 U2 ( .A1(n23), .A2(n24), .ZN(to_7[29]) );
  LVT_NAND2HSV8 U3 ( .A1(n47), .A2(n48), .ZN(to_7[17]) );
  LVT_INHSV4 U4 ( .I(n69), .ZN(n72) );
  LVT_CLKNHSV5 U5 ( .I(l_ctr), .ZN(n82) );
  LVT_INHSV0SR U6 ( .I(to_7[12]), .ZN(n2) );
  LVT_INHSV2 U7 ( .I(n2), .ZN(n14) );
  LVT_NAND2HSV8 U8 ( .A1(n27), .A2(n28), .ZN(to_7[7]) );
  LVT_CLKNAND2HSV8 U9 ( .A1(t_i_2_out[7]), .A2(n94), .ZN(n28) );
  LVT_CLKNAND2HSV3 U10 ( .A1(n59), .A2(n60), .ZN(to_7[13]) );
  LVT_NAND2HSV16 U11 ( .A1(n54), .A2(n55), .ZN(to_7[12]) );
  LVT_CLKNHSV12 U12 ( .I(n39), .ZN(n67) );
  LVT_IAO22HSV4 U13 ( .B1(t_i_2_out[0]), .B2(n94), .A1(n40), .A2(n94), .ZN(n39) );
  LVT_CLKNAND2HSV4 U14 ( .A1(n45), .A2(n46), .ZN(to_7[25]) );
  LVT_CLKNAND2HSV3 U15 ( .A1(t_i_2_out[25]), .A2(n94), .ZN(n46) );
  LVT_CLKNHSV12 U16 ( .I(n41), .ZN(n76) );
  LVT_IAO22HSV4 U17 ( .B1(t_i_2_out[3]), .B2(n94), .A1(n42), .A2(n94), .ZN(n41) );
  LVT_INHSV6 U18 ( .I(n63), .ZN(n73) );
  LVT_INHSV6SR U19 ( .I(n65), .ZN(n66) );
  LVT_CLKAND2HSV4 U20 ( .A1(t_i_2_out[28]), .A2(n94), .Z(n57) );
  LVT_NAND2HSV8 U21 ( .A1(t_i_2_out[12]), .A2(n94), .ZN(n55) );
  LVT_INHSV8 U22 ( .I(n29), .ZN(n30) );
  LVT_CLKNHSV3 U23 ( .I(mux_bq[31]), .ZN(n29) );
  LVT_INHSV2 U24 ( .I(n19), .ZN(n20) );
  LVT_INHSV2 U25 ( .I(l_g[24]), .ZN(n19) );
  LVT_CLKNHSV4 U26 ( .I(n64), .ZN(n74) );
  LVT_INHSV10 U27 ( .I(n31), .ZN(n32) );
  LVT_INHSV4SR U28 ( .I(n35), .ZN(n78) );
  LVT_MAOI22HSV4 U29 ( .A1(t_i_2_out[20]), .A2(n94), .B1(n36), .B2(n94), .ZN(
        n35) );
  LVT_INOR2HSV0 U30 ( .A1(l_t_i_1_in_0), .B1(n93), .ZN(c_t_i_1_in_0) );
  LVT_CLKNAND2HSV8 U31 ( .A1(n15), .A2(n16), .ZN(to_7[22]) );
  LVT_INHSV4 U32 ( .I(n53), .ZN(n15) );
  LVT_INHSV2 U33 ( .I(n52), .ZN(n16) );
  LVT_INHSV0SR U34 ( .I(to_7[2]), .ZN(n17) );
  LVT_INHSV2 U67 ( .I(n17), .ZN(n18) );
  LVT_INHSV4 U68 ( .I(n37), .ZN(n79) );
  LVT_INHSV4SR U70 ( .I(n68), .ZN(n70) );
  LVT_CLKNHSV5 U81 ( .I(l_g[27]), .ZN(n21) );
  LVT_INHSV10SR U82 ( .I(n21), .ZN(n22) );
  LVT_CLKNHSV5 U83 ( .I(n71), .ZN(n77) );
  LVT_AOI22HSV4 U84 ( .A1(ti_7[30]), .A2(ctro), .B1(t_i_2_out[30]), .B2(n94), 
        .ZN(n71) );
  LVT_CLKNHSV4 U85 ( .I(n51), .ZN(n75) );
  LVT_CLKNHSV6 U86 ( .I(to_7[6]), .ZN(n31) );
  LVT_CLKNAND2HSV2 U87 ( .A1(t_i_2_out[13]), .A2(n94), .ZN(n60) );
  LVT_CLKNAND2HSV4 U88 ( .A1(n43), .A2(n44), .ZN(to_7[21]) );
  LVT_CLKNAND2HSV8 U89 ( .A1(n80), .A2(n81), .ZN(to_1) );
  LVT_NAND2HSV3 U90 ( .A1(l_ctr), .A2(ti_1), .ZN(n80) );
  LVT_CLKNAND2HSV3 U91 ( .A1(t_i_2_out[21]), .A2(n94), .ZN(n44) );
  LVT_CLKNAND2HSV3 U92 ( .A1(t_i_2_out[29]), .A2(n94), .ZN(n24) );
  LVT_NAND2HSV4 U93 ( .A1(n49), .A2(n50), .ZN(to_7[8]) );
  LVT_OR2HSV16RD U94 ( .A1(n57), .A2(n56), .Z(to_7[28]) );
  LVT_AO22HSV4 U95 ( .A1(ti_7[23]), .A2(ctro), .B1(t_i_2_out[23]), .B2(n94), 
        .Z(to_7[23]) );
  LVT_MAOI22HSV2 U96 ( .A1(t_i_2_out[10]), .A2(n94), .B1(n38), .B2(n94), .ZN(
        n37) );
  LVT_CLKNAND2HSV2 U97 ( .A1(t_i_2_out[8]), .A2(n94), .ZN(n50) );
  LVT_NAND2HSV0 U98 ( .A1(ti_7[29]), .A2(ctro), .ZN(n23) );
  LVT_NAND2HSV16 U99 ( .A1(n25), .A2(n26), .ZN(to_7[1]) );
  LVT_CLKNAND2HSV8 U100 ( .A1(t_i_2_out[1]), .A2(n94), .ZN(n26) );
  LVT_CLKNAND2HSV8 U101 ( .A1(t_i_2_out[2]), .A2(n94), .ZN(n62) );
  LVT_NAND2HSV4 U102 ( .A1(t_i_2_out[17]), .A2(n94), .ZN(n48) );
  LVT_INHSV2 U103 ( .I(ti_7[10]), .ZN(n38) );
  LVT_INHSV2 U104 ( .I(ti_7[20]), .ZN(n36) );
  LVT_INHSV6 U105 ( .I(ctro), .ZN(n94) );
  LVT_INHSV2 U106 ( .I(ti_7[0]), .ZN(n40) );
  LVT_INHSV2 U107 ( .I(ti_7[3]), .ZN(n42) );
  LVT_NAND2HSV2 U108 ( .A1(ti_7[1]), .A2(ctro), .ZN(n25) );
  LVT_NAND2HSV2 U109 ( .A1(ti_7[7]), .A2(ctro), .ZN(n27) );
  LVT_AO22HSV4 U110 ( .A1(ti_7[15]), .A2(ctro), .B1(t_i_2_out[15]), .B2(n94), 
        .Z(n33) );
  LVT_INHSV2 U111 ( .I(n58), .ZN(n34) );
  LVT_NAND2HSV16 U112 ( .A1(n61), .A2(n62), .ZN(to_7[2]) );
  LVT_AND2HSV8 U113 ( .A1(t_i_2_out[22]), .A2(n94), .Z(n53) );
  LVT_NAND2HSV0 U114 ( .A1(ti_7[21]), .A2(ctro), .ZN(n43) );
  LVT_NAND2HSV0 U115 ( .A1(ti_7[25]), .A2(ctro), .ZN(n45) );
  LVT_NAND2HSV0 U116 ( .A1(ti_7[17]), .A2(ctro), .ZN(n47) );
  LVT_NAND2HSV0 U117 ( .A1(ti_7[8]), .A2(ctro), .ZN(n49) );
  LVT_INHSV0SR U118 ( .I(l_ctr), .ZN(n93) );
  LVT_CLKNAND2HSV8 U119 ( .A1(l_t_i_1_in_0), .A2(n82), .ZN(n81) );
  LVT_AOI22HSV4 U120 ( .A1(ti_7[5]), .A2(ctro), .B1(t_i_2_out[5]), .B2(n94), 
        .ZN(n51) );
  LVT_AND2HSV0RD U121 ( .A1(ti_7[22]), .A2(ctro), .Z(n52) );
  LVT_NAND2HSV0 U122 ( .A1(ti_7[12]), .A2(ctro), .ZN(n54) );
  LVT_AND2HSV0RD U123 ( .A1(ti_7[28]), .A2(ctro), .Z(n56) );
  LVT_INHSV2SR U124 ( .I(n93), .ZN(n58) );
  LVT_NAND2HSV0 U125 ( .A1(ti_7[13]), .A2(ctro), .ZN(n59) );
  LVT_NAND2HSV0 U126 ( .A1(ti_7[2]), .A2(ctro), .ZN(n61) );
  LVT_AOI22HSV4 U127 ( .A1(ti_7[19]), .A2(ctro), .B1(t_i_2_out[19]), .B2(n94), 
        .ZN(n63) );
  LVT_AOI22HSV4 U128 ( .A1(ti_7[18]), .A2(ctro), .B1(t_i_2_out[18]), .B2(n94), 
        .ZN(n64) );
  LVT_AOI22HSV4 U129 ( .A1(ti_7[26]), .A2(ctro), .B1(t_i_2_out[26]), .B2(n94), 
        .ZN(n65) );
  LVT_AOI22HSV4 U130 ( .A1(ti_7[9]), .A2(ctro), .B1(t_i_2_out[9]), .B2(n94), 
        .ZN(n68) );
  LVT_AOI22HSV4 U131 ( .A1(ti_7[27]), .A2(ctro), .B1(t_i_2_out[27]), .B2(n94), 
        .ZN(n69) );
  LVT_AO22HSV4 U132 ( .A1(ti_7[16]), .A2(ctro), .B1(t_i_2_out[16]), .B2(n94), 
        .Z(to_7[16]) );
  LVT_AO22HSV4 U133 ( .A1(ti_7[6]), .A2(ctro), .B1(t_i_2_out[6]), .B2(n94), 
        .Z(to_7[6]) );
  LVT_AO22HSV4 U134 ( .A1(ti_7[14]), .A2(ctro), .B1(t_i_2_out[14]), .B2(n94), 
        .Z(to_7[14]) );
  LVT_AO22HSV4 U135 ( .A1(ti_7[24]), .A2(ctro), .B1(t_i_2_out[24]), .B2(n94), 
        .Z(to_7[24]) );
  LVT_AO22HSV4 U136 ( .A1(ti_7[4]), .A2(ctro), .B1(t_i_2_out[4]), .B2(n94), 
        .Z(to_7[4]) );
  LVT_AO22HSV4 U137 ( .A1(ti_7[11]), .A2(ctro), .B1(t_i_2_out[11]), .B2(n94), 
        .Z(to_7[11]) );
endmodule


module regist_32bit_17 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV4 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV4 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV4 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV4 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n2), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n2), .Q(out[31]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n1), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n1), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n1), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n1), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n1), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n1), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n1), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n2), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n2), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n2), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_CLKNHSV4 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_32bit_16 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV2 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n2), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n2), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n2), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_32bit_15 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV4 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV4 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV4 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n2), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n2), .Q(out[31]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n1), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n1), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n1), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n1), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n1), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n2), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n2), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n2), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV4 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n1), .Q(out[19]) );
  LVT_DRNQHSV4 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV4 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n1), .Q(out[18]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_CLKNHSV4 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_1bit_11 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_10 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_31bit_11 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n1), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n1), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n1), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n1), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n1), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n1), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n1), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n2) );
  LVT_CLKNHSV4 U4 ( .I(n2), .ZN(n1) );
endmodule


module regist_31bit_10 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n1), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n2), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n2), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n1), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n2), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n2), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n1), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n2), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n2), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n2), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n2), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_INHSV2 U3 ( .I(n3), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n2) );
endmodule


module regist_1bit_9 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_32bit_14 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV4 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n2), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n2), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n2), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n2), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n2), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n2), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n2), .Q(out[27]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_CLKNHSV4 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_1bit_8 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_31bit_9 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n2), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n2), .Q(out[28]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n2), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n2), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n2), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n2), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n1) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n2) );
endmodule


module cell_3_2885 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_92 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_91 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_90 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_89 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_88 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_87 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_86 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_85 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_84 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_83 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_82 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_81 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_80 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_79 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_78 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_77 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_76 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_75 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_74 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_73 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV2 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_72 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_71 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_70 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_69 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_68 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U3 ( .A1(n5), .A2(n6), .Z(n7) );
endmodule


module cell_4_67 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV2 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n5), .A2(n6), .Z(n7) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_66 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n2), .A3(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_65 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_XOR3HSV1 U2 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
endmodule


module cell_4_64 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_63 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n2), .A3(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_62 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  LVT_NAND2HSV4 U1 ( .A1(n1), .A2(n3), .ZN(n6) );
  LVT_INHSV3SR U2 ( .I(n14), .ZN(n1) );
  LVT_CLKNAND2HSV2 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n13) );
  LVT_INHSV2 U4 ( .I(n13), .ZN(n8) );
  LVT_CLKNAND2HSV4 U5 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNAND2HSV0 U6 ( .A1(n12), .A2(n13), .ZN(n9) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n9), .A2(n10), .ZN(n14) );
  LVT_NAND2HSV2 U8 ( .A1(n11), .A2(n14), .ZN(n5) );
  LVT_CLKNAND2HSV3 U9 ( .A1(n8), .A2(n7), .ZN(n10) );
  LVT_INHSV1 U10 ( .I(n12), .ZN(n7) );
  LVT_XNOR2HSV1 U11 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n11) );
  LVT_AND2HSV2RD U12 ( .A1(b_in), .A2(a_in), .Z(n12) );
  LVT_INHSV2 U13 ( .I(n11), .ZN(n3) );
endmodule


module row_1_2 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [31:0] t_i_1_in;
  input [30:0] t_i_2_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_3_2885 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_92 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(t_i_1_out[1])
         );
  cell_4_91 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(t_i_1_out[2])
         );
  cell_4_90 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(t_i_1_out[3])
         );
  cell_4_89 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(t_i_1_out[4])
         );
  cell_4_88 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(t_i_1_out[5])
         );
  cell_4_87 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(t_i_1_out[6])
         );
  cell_4_86 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(t_i_1_out[7])
         );
  cell_4_85 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_2_in(t_i_2_in[7]), .t_i_out(t_i_1_out[8])
         );
  cell_4_84 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[9]), .t_i_2_in(t_i_2_in[8]), .t_i_out(t_i_1_out[9])
         );
  cell_4_83 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_2_in(t_i_2_in[9]), .t_i_out(
        t_i_1_out[10]) );
  cell_4_82 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[11]), .t_i_2_in(t_i_2_in[10]), .t_i_out(
        t_i_1_out[11]) );
  cell_4_81 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_2_in(t_i_2_in[11]), .t_i_out(
        t_i_1_out[12]) );
  cell_4_80 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_2_in(t_i_2_in[12]), .t_i_out(
        t_i_1_out[13]) );
  cell_4_79 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_2_in(t_i_2_in[13]), .t_i_out(
        t_i_1_out[14]) );
  cell_4_78 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_2_in(t_i_2_in[14]), .t_i_out(
        t_i_1_out[15]) );
  cell_4_77 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[16]), .t_i_2_in(t_i_2_in[15]), .t_i_out(
        t_i_1_out[16]) );
  cell_4_76 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_2_in(t_i_2_in[16]), .t_i_out(
        t_i_1_out[17]) );
  cell_4_75 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_2_in(t_i_2_in[17]), .t_i_out(
        t_i_1_out[18]) );
  cell_4_74 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_2_in(t_i_2_in[18]), .t_i_out(
        t_i_1_out[19]) );
  cell_4_73 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_2_in(t_i_2_in[19]), .t_i_out(
        t_i_1_out[20]) );
  cell_4_72 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_2_in(t_i_2_in[20]), .t_i_out(
        t_i_1_out[21]) );
  cell_4_71 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_2_in(t_i_2_in[21]), .t_i_out(
        t_i_1_out[22]) );
  cell_4_70 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_2_in(t_i_2_in[22]), .t_i_out(
        t_i_1_out[23]) );
  cell_4_69 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_2_in(t_i_2_in[23]), .t_i_out(
        t_i_1_out[24]) );
  cell_4_68 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_2_in(t_i_2_in[24]), .t_i_out(
        t_i_1_out[25]) );
  cell_4_67 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_2_in(t_i_2_in[25]), .t_i_out(
        t_i_1_out[26]) );
  cell_4_66 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_2_in(t_i_2_in[26]), .t_i_out(
        t_i_1_out[27]) );
  cell_4_65 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_2_in(t_i_2_in[27]), .t_i_out(
        t_i_1_out[28]) );
  cell_4_64 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_2_in(t_i_2_in[28]), .t_i_out(
        t_i_1_out[29]) );
  cell_4_63 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_2_in(t_i_2_in[29]), .t_i_out(
        t_i_1_out[30]) );
  cell_4_62 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[31]), .t_i_2_in(t_i_2_in[30]), .t_i_out(
        t_i_2_out) );
  LVT_BUFHSV2RT U1 ( .I(t_m_1_in), .Z(n1) );
  LVT_BUFHSV2RT U2 ( .I(t_m_1_in), .Z(n2) );
endmodule


module cell_2_92 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_2884 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2883 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2882 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2881 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2880 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2879 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2878 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2877 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2876 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2875 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2874 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2873 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2872 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2871 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2870 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2869 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2868 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2867 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2866 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2865 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2864 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2863 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2862 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2861 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2860 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2859 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2858 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2857 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2856 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2855 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2854 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV4 U1 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_CLKNAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV1 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2SR U5 ( .I(n7), .ZN(n4) );
  LVT_INHSV4SR U6 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_92 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_92 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2884 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2883 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2882 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2881 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2880 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2879 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2878 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2877 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2876 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2875 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2874 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2873 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2872 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2871 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2870 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2869 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2868 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2867 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2866 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2865 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2864 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2863 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2862 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2861 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2860 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2859 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2858 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2857 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2856 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2855 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2854 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV4SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV8 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_91 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_2853 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2852 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2851 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2850 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2849 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2848 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2847 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2846 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2845 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2844 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2843 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2842 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2841 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2840 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2839 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2838 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2837 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2836 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2835 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2834 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2833 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2832 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2831 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2830 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2829 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2828 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2827 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV1 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2826 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_INAND2HSV2 U1 ( .A1(n9), .B1(n8), .ZN(n6) );
  LVT_CLKNAND2HSV1 U2 ( .A1(n9), .A2(n4), .ZN(n5) );
  LVT_NAND2HSV2 U4 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNHSV2P5 U5 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XOR2HSV4 U7 ( .A1(n7), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_3_2825 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV4 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV3SR U5 ( .I(n9), .ZN(n2) );
  LVT_INHSV2SR U6 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV0P5 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV1 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module cell_3_2824 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_CLKNHSV0P5 U1 ( .I(n8), .ZN(n2) );
  LVT_IOA21HSV4 U2 ( .A1(n2), .A2(n4), .B(n5), .ZN(t_i_out) );
  LVT_CLKNHSV2 U4 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0P5 U5 ( .A1(n8), .A2(n6), .ZN(n5) );
  LVT_NAND2HSV0P5 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XNOR2HSV4 U7 ( .A1(t_i_1_in), .A2(n7), .ZN(n6) );
endmodule


module cell_3_2823 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV1 U1 ( .A1(n5), .A2(n9), .ZN(n7) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_NAND2HSV2 U3 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(n10), .A2(n4), .ZN(n6) );
  LVT_CLKNHSV2 U5 ( .I(n10), .ZN(n5) );
  LVT_NAND2HSV2 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_XNOR2HSV4 U7 ( .A1(n8), .A2(t_i_1_in), .ZN(n4) );
  LVT_NAND2HSV0 U8 ( .A1(b_in), .A2(a_in), .ZN(n8) );
endmodule


module row_other_91 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1;

  cell_2_91 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2853 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2852 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2851 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2850 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2849 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2848 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2847 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2846 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2845 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2844 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2843 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2842 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2841 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2840 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2839 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2838 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2837 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2836 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2835 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2834 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2833 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2832 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2831 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2830 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2829 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2828 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2827 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2826 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2825 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2824 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2823 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV6RQ U1 ( .I(t_m_1_in), .Z(n1) );
endmodule


module cell_2_90 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_2822 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2821 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2820 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2819 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2818 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2817 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2816 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2815 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2814 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2813 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2812 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2811 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2810 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2809 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2808 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2807 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2806 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2805 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2804 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2803 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2802 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2801 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2800 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2799 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2798 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2797 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2796 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2795 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_2794 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2793 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_2792 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV3SR U1 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV3 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNHSV2P5 U5 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_90 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_90 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2822 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2821 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2820 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2819 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2818 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2817 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2816 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2815 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2814 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2813 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2812 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2811 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2810 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2809 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2808 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2807 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2806 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2805 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2804 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2803 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2802 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2801 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2800 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2799 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2798 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2797 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2796 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2795 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2794 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2793 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2792 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV6 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_89 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_2791 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2790 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2789 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2788 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2787 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2786 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2785 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2784 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2783 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2782 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2781 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2780 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2779 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2778 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2777 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2776 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2775 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2774 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2773 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2772 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2771 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2770 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2769 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2768 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2767 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XOR2HSV0 U4 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_2766 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2765 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2764 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2763 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2762 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_2761 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4, n5;

  LVT_NAND2HSV0P5 U1 ( .A1(n5), .A2(n4), .ZN(n3) );
  LVT_CLKXOR2HSV2 U2 ( .A1(t_i_1_in), .A2(n2), .Z(n4) );
  LVT_OAI21HSV2 U3 ( .A1(n4), .A2(n5), .B(n3), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKAND2HSV2 U5 ( .A1(b_in), .A2(a_in), .Z(n2) );
endmodule


module row_other_89 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_89 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2791 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2790 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2789 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2788 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2787 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2786 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2785 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2784 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2783 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2782 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2781 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2780 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2779 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2778 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2777 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2776 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2775 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2774 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2773 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2772 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2771 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2770 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2769 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2768 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2767 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2766 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2765 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2764 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2763 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2762 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2761 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV4 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV2 U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_88 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_2760 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2759 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2758 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2757 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2756 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2755 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2754 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2753 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2752 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2751 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2750 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2749 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2748 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2747 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2746 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2745 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2744 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2743 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2742 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2741 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2740 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2739 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2738 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2737 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2736 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2735 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2734 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2733 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2732 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2731 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2730 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_88 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_88 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2760 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2759 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2758 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2757 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2756 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2755 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2754 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2753 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2752 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2751 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2750 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2749 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2748 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2747 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2746 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2745 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2744 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2743 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2742 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2741 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2740 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2739 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2738 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2737 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2736 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2735 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2734 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2733 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2732 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2731 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2730 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2 U1 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n2), .ZN(n3) );
  LVT_INHSV0SR U3 ( .I(t_m_1_in), .ZN(n2) );
endmodule


module cell_2_87 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_2729 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2728 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2727 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2726 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2725 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2724 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2723 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2722 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2721 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2720 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2719 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2718 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2717 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2716 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2715 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2714 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2713 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2712 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2711 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2710 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2709 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2708 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2707 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2706 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2705 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2704 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2703 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2702 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2701 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2700 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2699 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module row_other_87 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4, n5, n6;

  cell_2_87 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2729 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2728 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2727 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2726 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2725 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2724 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2723 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2722 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2721 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2720 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2719 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2718 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2717 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2716 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2715 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2714 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2713 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2712 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2711 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2710 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2709 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2708 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2707 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2706 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2705 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2704 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2703 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2702 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2701 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2700 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2699 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV10 U1 ( .I(n1), .ZN(n3) );
  LVT_INHSV8SR U2 ( .I(n6), .ZN(n1) );
  LVT_INHSV4SR U3 ( .I(n4), .ZN(n6) );
  LVT_INHSV4 U4 ( .I(t_m_1_in), .ZN(n4) );
  LVT_INHSV1SR U5 ( .I(n1), .ZN(n2) );
  LVT_INHSV2 U6 ( .I(n4), .ZN(n5) );
endmodule


module cell_2_86 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_2698 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2697 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2696 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2695 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2694 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2693 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2692 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2691 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2690 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2689 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2688 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2687 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2686 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2685 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2684 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2683 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2682 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2681 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2680 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2679 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2678 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2677 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2676 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2675 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2674 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2673 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2672 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2671 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2670 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2669 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2668 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module row_other_86 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_86 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2698 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2697 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2696 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2695 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2694 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2693 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2692 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2691 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2690 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2689 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2688 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2687 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2686 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2685 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2684 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2683 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2682 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2681 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2680 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2679 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2678 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2677 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2676 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2675 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2674 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2673 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2672 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2671 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2670 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2669 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2668 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV4 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_85 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_2667 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2666 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2665 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2664 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2663 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2662 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2661 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2660 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2659 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2658 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2657 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2656 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2655 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2654 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2653 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2652 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2651 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2650 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2649 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2648 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2647 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2646 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2645 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2644 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV4 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2643 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2642 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2641 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2640 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2639 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2638 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2637 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(g_in), .A2(t_m_1_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_85 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_85 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2667 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2666 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2665 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2664 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2663 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2662 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2661 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2660 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2659 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2658 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2657 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2656 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2655 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2654 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2653 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2652 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2651 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2650 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2649 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2648 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2647 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2646 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2645 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2644 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2643 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2642 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2641 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2640 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2639 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2638 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2637 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV0P5SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV6SR U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_84 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_2636 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2635 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2634 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2633 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2632 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2631 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2630 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2629 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2628 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2627 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2626 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2625 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2624 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2623 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2622 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2621 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2620 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2619 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2618 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2617 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2616 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2615 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2614 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2613 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2612 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2611 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2610 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2609 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2608 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2607 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2606 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV2P5 U1 ( .I(n7), .ZN(n4) );
  LVT_INHSV3SR U2 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV1 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV4 U5 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV4 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_84 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4, n5;

  cell_2_84 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2636 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2635 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2634 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2633 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2632 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2631 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2630 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2629 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2628 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2627 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2626 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2625 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2624 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2623 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2622 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2621 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2620 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2619 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2618 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2617 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2616 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2615 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2614 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2613 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2612 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2611 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2610 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2609 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2608 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2607 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2606 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV8 U1 ( .I(n1), .ZN(n3) );
  LVT_INHSV4 U2 ( .I(n4), .ZN(n1) );
  LVT_INHSV2SR U3 ( .I(n5), .ZN(n4) );
  LVT_INHSV2SR U4 ( .I(t_m_1_in), .ZN(n5) );
  LVT_INHSV0P5 U5 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_83 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_2605 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2604 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2603 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2602 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2601 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2600 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2599 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2598 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2597 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2596 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2595 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2594 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2593 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2592 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2591 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2590 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2589 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2588 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2587 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2586 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2585 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2584 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2583 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2582 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2581 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2580 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV2 U1 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_OR2HSV1RD U2 ( .A1(n4), .A2(t_i_1_in), .Z(n6) );
  LVT_INHSV2 U3 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0P5 U5 ( .A1(n5), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U6 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_CLKNHSV0P5 U7 ( .I(n8), .ZN(n5) );
  LVT_XOR2HSV2 U8 ( .A1(n10), .A2(n9), .Z(t_i_out) );
endmodule


module cell_3_2579 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2578 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2577 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2576 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2575 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV2SR U1 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV3 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV2 U4 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV2SR U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV1 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_XNOR2HSV1 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_83 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_83 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_2605 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2604 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2603 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2602 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2601 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2600 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2599 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2598 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2597 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2596 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2595 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2594 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2593 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2592 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2591 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2590 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2589 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2588 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2587 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2586 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2585 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2584 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2583 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2582 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2581 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2580 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2579 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2578 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2577 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2576 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2575 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_82 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_2574 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2573 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2572 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2571 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2570 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2569 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2568 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2567 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2566 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2565 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2564 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2563 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2562 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2561 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2560 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2559 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2558 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2557 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2556 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2555 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2554 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2553 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2552 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2551 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2550 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2549 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_NAND2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U5 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV1 U6 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_3_2548 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2547 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2546 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2545 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_2544 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XNOR2HSV4 U1 ( .A1(n8), .A2(t_i_1_in), .ZN(n4) );
  LVT_NAND2HSV1 U2 ( .A1(n9), .A2(n4), .ZN(n6) );
  LVT_INHSV2SR U4 ( .I(n9), .ZN(n5) );
  LVT_CLKNAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV2 U6 ( .A1(n7), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U7 ( .A1(n5), .A2(n2), .ZN(n7) );
  LVT_XOR2HSV0 U8 ( .A1(n8), .A2(t_i_1_in), .Z(n2) );
endmodule


module row_other_82 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_82 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2574 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2573 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2572 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2571 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2570 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2569 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2568 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2567 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2566 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2565 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2564 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2563 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2562 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2561 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2560 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2559 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2558 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2557 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2556 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2555 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2554 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2553 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2552 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2551 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2550 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2549 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2548 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2547 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2546 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2545 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2544 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV4RT U1 ( .I(n2), .Z(n1) );
  LVT_BUFHSV6RQ U2 ( .I(t_m_1_in), .Z(n2) );
endmodule


module cell_2_81 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_2543 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2542 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2541 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2540 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2539 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2538 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2537 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2536 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2535 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2534 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2533 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2532 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2531 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2530 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2529 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2528 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2527 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2526 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2525 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2524 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2523 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2522 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2521 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2520 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2519 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2518 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U3 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_2517 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2516 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2515 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2514 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_INHSV2SR U1 ( .I(n8), .ZN(n4) );
  LVT_OAI21HSV2 U4 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_NAND2HSV2 U6 ( .A1(n4), .A2(n7), .ZN(n5) );
endmodule


module cell_3_2513 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV1 U1 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV3 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV2 U4 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNHSV2P5 U5 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV3SR U7 ( .I(n9), .ZN(n2) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_81 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_81 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2543 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2542 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2541 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2540 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2539 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2538 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2537 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2536 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2535 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2534 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2533 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2532 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2531 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2530 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2529 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2528 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2527 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2526 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2525 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2524 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2523 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2522 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2521 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2520 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2519 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2518 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2517 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2516 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2515 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2514 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2513 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV3SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV10 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_80 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_2512 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2511 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2510 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2509 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2508 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2507 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2506 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2505 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2504 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2503 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2502 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2501 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2500 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2499 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2498 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2497 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2496 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2495 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2494 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2493 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2492 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2491 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV0P5 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_2490 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2489 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2488 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2487 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2486 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2485 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2484 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XOR2HSV2 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0P5 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_2483 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_CLKNHSV0P5 U4 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XOR2HSV4 U6 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
endmodule


module cell_3_2482 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module row_other_80 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_2_80 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2512 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2511 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2510 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2509 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2508 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2507 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2506 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2505 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2504 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2503 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2502 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2501 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2500 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2499 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2498 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2497 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2496 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2495 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2494 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2493 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2492 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2491 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2490 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2489 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2488 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2487 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2486 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2485 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2484 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2483 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2482 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2SR U1 ( .I(t_m_1_in), .ZN(n3) );
  LVT_CLKNHSV4 U2 ( .I(n3), .ZN(n4) );
  LVT_CLKNHSV2 U3 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U4 ( .I(n4), .ZN(n1) );
endmodule


module cell_2_79 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_2481 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2480 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2479 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2478 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2477 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2476 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2475 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2474 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2473 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2472 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2471 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2470 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2469 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2468 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2467 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2466 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2465 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2464 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2463 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2462 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2461 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2460 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2459 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2458 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2457 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2456 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2455 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2454 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2453 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV0 U4 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U5 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_2452 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV3 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV1 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNAND2HSV3 U3 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0SR U4 ( .I(n8), .ZN(n4) );
  LVT_INHSV2P5 U5 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV0 U6 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV2 U7 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_2451 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV4 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module row_other_79 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_79 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2481 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2480 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2479 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2478 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2477 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2476 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2475 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2474 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2473 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2472 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2471 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2470 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2469 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2468 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2467 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2466 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2465 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2464 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2463 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2462 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2461 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2460 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2459 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2458 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2457 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2456 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2455 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2454 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2453 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2452 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2451 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV16SR U1 ( .I(n1), .ZN(n2) );
  LVT_CLKNHSV12 U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_78 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_2450 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2449 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2448 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2447 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2446 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2445 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2444 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2443 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2442 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2441 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2440 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2439 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2438 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2437 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2436 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2435 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2434 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2433 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2432 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2431 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2430 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2429 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2428 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2427 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2426 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2425 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2424 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2423 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2422 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2421 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2420 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U4 ( .I(n7), .ZN(n4) );
  LVT_INHSV3SR U5 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV2 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV0P5 U7 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_78 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_78 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2450 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2449 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2448 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2447 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2446 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2445 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2444 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2443 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2442 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2441 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2440 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2439 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2438 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2437 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2436 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2435 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2434 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2433 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2432 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2431 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2430 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2429 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2428 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2427 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2426 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2425 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2424 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2423 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2422 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2421 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2420 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV1SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_77 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_2419 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2418 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2417 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2416 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2415 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2414 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2413 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2412 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2411 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2410 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2409 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2408 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2407 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2406 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2405 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2404 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2403 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2402 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2401 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2400 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2399 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2398 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2397 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2396 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2395 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2394 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2393 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2392 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2391 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2390 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11;

  LVT_NAND2HSV4 U1 ( .A1(n4), .A2(n5), .ZN(n9) );
  LVT_NAND2HSV1 U2 ( .A1(n10), .A2(t_i_1_in), .ZN(n4) );
  LVT_CLKNAND2HSV3 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n11) );
  LVT_INHSV3SR U4 ( .I(n11), .ZN(n6) );
  LVT_NOR2HSV2 U5 ( .A1(n10), .A2(t_i_1_in), .ZN(n2) );
  LVT_INHSV2SR U6 ( .I(n2), .ZN(n5) );
  LVT_IOA21HSV4 U7 ( .A1(n11), .A2(n9), .B(n8), .ZN(t_i_out) );
  LVT_NAND2HSV0 U8 ( .A1(b_in), .A2(a_in), .ZN(n10) );
  LVT_INHSV3SR U9 ( .I(n9), .ZN(n7) );
  LVT_NAND2HSV4 U10 ( .A1(n6), .A2(n7), .ZN(n8) );
endmodule


module cell_3_2389 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV3 U1 ( .I(n9), .ZN(n2) );
  LVT_XNOR2HSV4 U2 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNHSV2 U4 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV4 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U7 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV3 U8 ( .A1(n2), .A2(n4), .ZN(n6) );
endmodule


module row_other_77 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_77 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2419 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2418 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2417 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2416 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2415 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2414 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2413 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2412 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2411 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2410 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2409 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2408 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2407 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2406 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2405 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2404 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2403 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2402 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2401 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2400 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2399 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2398 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2397 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2396 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2395 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2394 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2393 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2392 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2391 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2390 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2389 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2SR U1 ( .I(t_m_1_in), .ZN(n3) );
  LVT_INHSV2 U2 ( .I(n3), .ZN(n1) );
  LVT_INHSV2 U3 ( .I(n3), .ZN(n2) );
endmodule


module cell_2_76 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_2388 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2387 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2386 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2385 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2384 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2383 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2382 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2381 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2380 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2379 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2378 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2377 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2376 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2375 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2374 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2373 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2372 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2371 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2370 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2369 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2368 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2367 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2366 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2365 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_NAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV0 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_2364 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2363 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2362 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2361 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2360 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2359 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2358 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n8), .A2(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV2 U4 ( .A1(n5), .A2(n6), .ZN(n7) );
  LVT_INHSV2 U5 ( .I(n8), .ZN(n2) );
  LVT_INHSV2 U6 ( .I(t_i_1_in), .ZN(n4) );
  LVT_XNOR2HSV4 U7 ( .A1(n9), .A2(n7), .ZN(t_i_out) );
  LVT_NAND2HSV2 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
endmodule


module row_other_76 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_76 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2388 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2387 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2386 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2385 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2384 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2383 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2382 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2381 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2380 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2379 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2378 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2377 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2376 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2375 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2374 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2373 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2372 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2371 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2370 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2369 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2368 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2367 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2366 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2365 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2364 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2363 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2362 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2361 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2360 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2359 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2358 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_CLKNHSV12 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_75 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_2357 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2356 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2355 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2354 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2353 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2352 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2351 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2350 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2349 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2348 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2347 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2346 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2345 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2344 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2343 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2342 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2341 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2340 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2339 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2338 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2337 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2336 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2335 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2334 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2333 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2332 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2331 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2330 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2329 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_2328 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U3 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV0 U4 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U5 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U6 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_3_2327 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV4 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNHSV2 U2 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV0P5 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2 U5 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U6 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV4 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV4 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
endmodule


module row_other_75 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1;

  cell_2_75 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_2357 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2356 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2355 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2354 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2353 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2352 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2351 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2350 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2349 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2348 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2347 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2346 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2345 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2344 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2343 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2342 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2341 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2340 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2339 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2338 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2337 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2336 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2335 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2334 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2333 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2332 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2331 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2330 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2329 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2328 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2327 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV2RT U1 ( .I(t_m_1_in), .Z(n1) );
endmodule


module cell_2_74 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_2326 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2325 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2324 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2323 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2322 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2321 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2320 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2319 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2318 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2317 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2316 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2315 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2314 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2313 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2312 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2311 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2310 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2309 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2308 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2307 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2306 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2305 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2304 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2303 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV0P5 U5 ( .I(n6), .ZN(n4) );
  LVT_CLKNAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_2302 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2301 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2300 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
endmodule


module cell_3_2299 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV0 U2 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_CLKNAND2HSV2 U4 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_NAND2HSV2 U5 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_CLKNHSV2 U6 ( .I(n10), .ZN(n4) );
  LVT_INHSV0SR U7 ( .I(n9), .ZN(n5) );
  LVT_CLKXOR2HSV2 U8 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
endmodule


module cell_3_2298 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2297 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2296 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_NOR2HSV3 U1 ( .A1(n8), .A2(n6), .ZN(n2) );
  LVT_NAND2HSV2 U2 ( .A1(n4), .A2(n5), .ZN(t_i_out) );
  LVT_INHSV2SR U4 ( .I(n2), .ZN(n5) );
  LVT_XNOR2HSV4 U5 ( .A1(t_i_1_in), .A2(n7), .ZN(n6) );
  LVT_NAND2HSV0 U6 ( .A1(n8), .A2(n6), .ZN(n4) );
  LVT_NAND2HSV4 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module row_other_74 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_74 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2326 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2325 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2324 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2323 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2322 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2321 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2320 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2319 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2318 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2317 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2316 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2315 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2314 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2313 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2312 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2311 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2310 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2309 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2308 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2307 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2306 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2305 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2304 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2303 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2302 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2301 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2300 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2299 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2298 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2297 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2296 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV8 U1 ( .I(n1), .ZN(n2) );
  LVT_CLKNHSV4 U2 ( .I(n3), .ZN(n1) );
  LVT_BUFHSV2RT U3 ( .I(t_m_1_in), .Z(n3) );
endmodule


module cell_2_73 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_2295 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2294 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2293 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2292 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2291 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2290 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2289 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2288 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2287 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2286 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2285 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2284 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2283 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2282 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2281 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2280 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2279 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2278 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2277 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2276 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2275 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2274 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2273 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2272 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2271 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2270 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2269 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_XOR2HSV2 U1 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0P5SR U3 ( .I(n4), .ZN(n6) );
  LVT_INOR2HSV1 U5 ( .A1(n8), .B1(t_i_1_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U6 ( .A1(n5), .A2(t_i_1_in), .ZN(n7) );
  LVT_INHSV0SR U7 ( .I(n8), .ZN(n5) );
  LVT_NAND2HSV0 U8 ( .A1(b_in), .A2(a_in), .ZN(n8) );
endmodule


module cell_3_2268 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_NAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV1 U3 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV0P5 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_2267 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKXOR2HSV4 U2 ( .A1(n5), .A2(n6), .Z(t_i_out) );
endmodule


module cell_3_2266 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2265 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV4 U1 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV2 U5 ( .I(n9), .ZN(n2) );
  LVT_INHSV3 U6 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV1 U7 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_73 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1;

  cell_2_73 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2295 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2294 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2293 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2292 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2291 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2290 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2289 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2288 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2287 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2286 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2285 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2284 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2283 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2282 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2281 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2280 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2279 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2278 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2277 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2276 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2275 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2274 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2273 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2272 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2271 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2270 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2269 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2268 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2267 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2266 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2265 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV4 U1 ( .I(t_m_1_in), .Z(n1) );
endmodule


module cell_2_72 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_2264 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2263 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2262 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2261 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2260 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2259 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2258 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2257 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2256 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2255 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2254 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2253 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2252 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2251 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2250 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2249 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2248 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2247 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2246 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2245 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2244 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2243 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2242 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2241 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2240 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2239 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2238 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2237 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2236 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_2235 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV1 U1 ( .A1(n8), .A2(t_i_1_in), .Z(n2) );
  LVT_XNOR2HSV2 U2 ( .A1(n8), .A2(t_i_1_in), .ZN(n4) );
  LVT_INHSV2 U4 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV2 U5 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_NAND2HSV2 U6 ( .A1(n9), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV2 U7 ( .A1(n5), .A2(n2), .ZN(n7) );
  LVT_NAND2HSV2 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
endmodule


module cell_3_2234 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV1 U4 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2SR U5 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV0 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2 U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_72 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_72 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2264 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2263 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2262 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2261 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2260 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2259 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2258 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2257 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2256 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2255 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2254 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2253 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2252 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2251 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2250 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2249 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2248 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2247 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2246 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2245 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2244 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2243 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2242 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2241 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2240 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2239 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2238 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2237 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2236 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2235 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2234 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV6RT U1 ( .I(t_m_1_in), .Z(n2) );
  LVT_BUFHSV4RQ U2 ( .I(n2), .Z(n1) );
endmodule


module cell_2_71 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_2233 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2232 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2231 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2230 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2229 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2228 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2227 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2226 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2225 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2224 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2223 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2222 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2221 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2220 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2219 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2218 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2217 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2216 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2215 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2214 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2213 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2212 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2211 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2210 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2209 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2208 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2207 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2206 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2205 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2204 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U1 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV4 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV2SR U5 ( .I(n10), .ZN(n4) );
  LVT_CLKNHSV1 U6 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV0P5 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_XOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
endmodule


module cell_3_2203 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_71 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_71 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_2233 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2232 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2231 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2230 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2229 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2228 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2227 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2226 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2225 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2224 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2223 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2222 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2221 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2220 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2219 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2218 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2217 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2216 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2215 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2214 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2213 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2212 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2211 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2210 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2209 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2208 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2207 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2206 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2205 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2204 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2203 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_70 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_2202 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2201 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2200 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2199 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2198 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2197 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2196 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2195 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2194 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2193 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2192 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2191 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2190 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2189 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2188 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2187 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2186 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2185 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2184 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2183 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2182 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2181 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2180 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2179 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2178 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2177 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2176 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2175 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2174 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV1 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV0 U5 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_2173 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2172 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module row_other_70 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_70 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2202 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2201 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2200 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2199 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2198 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2197 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2196 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2195 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2194 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2193 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2192 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2191 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2190 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2189 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2188 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2187 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2186 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2185 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2184 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2183 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2182 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2181 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2180 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2179 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2178 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2177 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2176 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2175 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2174 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2173 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2172 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2 U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV8 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_69 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_2171 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2170 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2169 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2168 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2167 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2166 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2165 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2164 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2163 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2162 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2161 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2160 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2159 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2158 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2157 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2156 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2155 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2154 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2153 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2152 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2151 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2150 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2149 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2148 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2147 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2146 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2145 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2144 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XOR2HSV0 U4 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_2143 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2142 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2141 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n6), .B(n2), .ZN(t_i_out) );
  LVT_NAND2HSV4 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKNAND2HSV1 U4 ( .A1(n6), .A2(n4), .ZN(n2) );
  LVT_XNOR2HSV1 U5 ( .A1(n5), .A2(t_i_1_in), .ZN(n4) );
endmodule


module row_other_69 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_69 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2171 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2170 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2169 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2168 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2167 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2166 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2165 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2164 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2163 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2162 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2161 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2160 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2159 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2158 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2157 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2156 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2155 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2154 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2153 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2152 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2151 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2150 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2149 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2148 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2147 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2146 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2145 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2144 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2143 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2142 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2141 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV4 U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV8 U2 ( .I(n1), .ZN(n3) );
  LVT_INHSV4SR U3 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_68 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_2140 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2139 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2138 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2137 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2136 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2135 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2134 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2133 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2132 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2131 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2130 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2129 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2128 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2127 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2126 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2125 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2124 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2123 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2122 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2121 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2120 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2119 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2118 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2117 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2116 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2115 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2114 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2113 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2112 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2111 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n14) );
  LVT_CLKNAND2HSV0 U2 ( .A1(n4), .A2(n13), .ZN(n7) );
  LVT_CLKNAND2HSV1 U3 ( .A1(n10), .A2(n11), .ZN(n13) );
  LVT_INHSV2 U4 ( .I(n14), .ZN(n4) );
  LVT_NAND2HSV0P5 U5 ( .A1(n5), .A2(n14), .ZN(n6) );
  LVT_INHSV0SR U6 ( .I(n13), .ZN(n5) );
  LVT_NAND2HSV2 U7 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_NAND2HSV2 U8 ( .A1(n12), .A2(n9), .ZN(n10) );
  LVT_NAND2HSV2 U9 ( .A1(n8), .A2(t_i_1_in), .ZN(n11) );
  LVT_CLKNHSV0 U10 ( .I(n12), .ZN(n8) );
  LVT_INHSV2 U11 ( .I(t_i_1_in), .ZN(n9) );
  LVT_NAND2HSV0 U12 ( .A1(b_in), .A2(a_in), .ZN(n12) );
endmodule


module cell_3_2110 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_CLKNAND2HSV1 U1 ( .A1(n5), .A2(t_i_1_in), .ZN(n2) );
  LVT_OAI21HSV2 U2 ( .A1(t_i_1_in), .A2(n5), .B(n2), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XNOR2HSV4 U5 ( .A1(n4), .A2(n6), .ZN(t_i_out) );
endmodule


module row_other_68 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4, n5, n6, n7;

  cell_2_68 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2140 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2139 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2138 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2137 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2136 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2135 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2134 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2133 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2132 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2131 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2130 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2129 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n6), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2128 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2127 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2126 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2125 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n6), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2124 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2123 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2122 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2121 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2120 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2119 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2118 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2117 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2116 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2115 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n6), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2114 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n6), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2113 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2112 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2111 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        n5), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2110 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV2RT U1 ( .I(n4), .Z(n1) );
  LVT_BUFHSV8 U2 ( .I(n4), .Z(n2) );
  LVT_BUFHSV8 U3 ( .I(n4), .Z(n3) );
  LVT_CLKNHSV2P5 U4 ( .I(n7), .ZN(n4) );
  LVT_INHSV1SR U5 ( .I(n7), .ZN(n6) );
  LVT_INHSV4SR U6 ( .I(n7), .ZN(n5) );
  LVT_INHSV2SR U7 ( .I(t_m_1_in), .ZN(n7) );
endmodule


module cell_2_67 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_2109 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2108 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2107 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2106 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2105 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2104 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2103 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2102 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2101 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2100 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2099 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2098 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2097 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2096 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2095 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2094 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2093 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2092 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2091 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2090 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2089 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2088 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2087 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2086 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2085 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2084 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2083 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2082 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2081 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2080 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_INHSV2 U2 ( .I(n9), .ZN(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_NAND2HSV0P5 U5 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV2SR U7 ( .I(n10), .ZN(n4) );
  LVT_NAND2HSV0P5 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_2079 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_67 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_67 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2109 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2108 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2107 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2106 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2105 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2104 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2103 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2102 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2101 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2100 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2099 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2098 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2097 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2096 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2095 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2094 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2093 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2092 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2091 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2090 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2089 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2088 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2087 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2086 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2085 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2084 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2083 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2082 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2081 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2080 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2079 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV6 U1 ( .I(n2), .ZN(n3) );
  LVT_CLKNHSV2 U2 ( .I(t_m_1_in), .ZN(n2) );
  LVT_INHSV0P5SR U3 ( .I(n2), .ZN(n1) );
endmodule


module cell_2_66 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_2078 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2077 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2076 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2075 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2074 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2073 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2072 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2071 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2070 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2069 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2068 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2067 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2066 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2065 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2064 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2063 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2062 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2061 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2060 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2059 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2058 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2057 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2056 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2055 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2054 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2053 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2052 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2051 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U3 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV8 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKXOR2HSV2 U6 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_3_2050 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2049 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n2), .A2(n5), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_2048 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_66 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_66 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_2078 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2077 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2076 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2075 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2074 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2073 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2072 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2071 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2070 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2069 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2068 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2067 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2066 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2065 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2064 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2063 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2062 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2061 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2060 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2059 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2058 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2057 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2056 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2055 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2054 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2053 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2052 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2051 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2050 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2049 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2048 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV3 U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_CLKNHSV12 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_65 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_2047 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2046 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2045 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2044 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2043 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2042 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2041 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2040 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2039 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2038 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2037 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2036 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2035 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2034 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2033 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2032 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2031 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2030 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2029 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2028 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2027 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2026 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2025 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2024 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2023 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2022 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2021 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2020 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2019 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_2018 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2017 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_65 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_65 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_2047 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2046 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2045 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2044 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2043 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2042 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2041 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2040 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2039 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2038 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2037 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2036 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2035 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2034 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2033 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2032 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2031 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_2030 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_2029 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_2028 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_2027 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_2026 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_2025 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_2024 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_2023 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_2022 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_2021 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_2020 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2019 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_2018 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_2017 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV2 U1 ( .I(t_m_1_in), .ZN(n2) );
  LVT_INHSV6 U2 ( .I(n2), .ZN(n3) );
  LVT_CLKNHSV1 U3 ( .I(n2), .ZN(n1) );
endmodule


module cell_2_64 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_2016 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2015 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2014 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2013 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2012 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2011 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2010 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2009 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2008 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2007 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV2 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U5 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0SR U6 ( .I(n8), .ZN(n4) );
  LVT_INHSV2 U7 ( .I(t_i_1_in), .ZN(n5) );
  LVT_CLKXOR2HSV2 U8 ( .A1(n10), .A2(n9), .Z(t_i_out) );
endmodule


module cell_3_2006 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_2005 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2004 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2003 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2002 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2001 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_2000 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1999 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1998 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1997 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1996 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1995 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1994 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1993 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1992 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1991 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1990 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1989 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1988 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1987 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV1 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module cell_3_1986 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_CLKNAND2HSV2 U1 ( .A1(n6), .A2(n4), .ZN(n2) );
  LVT_OAI21HSV2 U2 ( .A1(n6), .A2(n4), .B(n2), .ZN(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XNOR2HSV4 U5 ( .A1(t_i_1_in), .A2(n5), .ZN(n4) );
endmodule


module row_other_64 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_64 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_2016 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_2015 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_2014 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_2013 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_2012 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_2011 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_2010 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_2009 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_2008 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_2007 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_2006 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_2005 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_2004 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_2003 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_2002 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_2001 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_2000 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1999 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1998 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1997 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1996 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1995 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1994 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1993 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1992 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1991 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1990 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1989 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1988 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1987 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1986 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV8 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV2 U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_63 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1985 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1984 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1983 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1982 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1981 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1980 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1979 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1978 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1977 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1976 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1975 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1974 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_XOR2HSV0 U1 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_CLKNAND2HSV2 U2 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_CLKNAND2HSV1 U3 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U5 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0SR U6 ( .I(n8), .ZN(n4) );
  LVT_CLKNHSV2P5 U7 ( .I(t_i_1_in), .ZN(n5) );
  LVT_CLKNAND2HSV8 U8 ( .A1(b_in), .A2(a_in), .ZN(n8) );
endmodule


module cell_3_1973 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1972 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1971 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1970 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1969 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV1 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_INHSV0SR U4 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XOR2HSV4 U6 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
endmodule


module cell_3_1968 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1967 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1966 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1965 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1964 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1963 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1962 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1961 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1960 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1959 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1958 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
endmodule


module cell_3_1957 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1956 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1955 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_CLKNAND2HSV3 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module row_other_63 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_63 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_1985 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1984 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1983 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1982 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1981 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1980 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1979 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1978 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1977 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1976 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1975 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1974 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1973 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1972 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1971 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1970 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1969 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1968 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1967 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1966 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1965 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1964 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1963 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1962 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1961 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1960 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1959 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1958 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1957 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1956 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1955 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_62 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_1954 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV0 U1 ( .A1(n4), .A2(n8), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(n8), .A2(n4), .ZN(n5) );
  LVT_INHSV0SR U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_1953 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV0 U1 ( .A1(n4), .A2(n8), .B(n5), .ZN(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U4 ( .A1(n8), .A2(n4), .ZN(n5) );
  LVT_INHSV0SR U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_1952 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_INHSV2SR U2 ( .I(n8), .ZN(n4) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_1951 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_INHSV2SR U2 ( .I(n8), .ZN(n4) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_1950 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_INHSV2SR U2 ( .I(n8), .ZN(n4) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_1949 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_INHSV2SR U2 ( .I(n8), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(g_in), .A2(t_m_1_in), .ZN(n8) );
  LVT_XOR2HSV0 U5 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U6 ( .A1(n4), .A2(n7), .ZN(n5) );
endmodule


module cell_3_1948 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_INHSV2SR U2 ( .I(n8), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(g_in), .A2(t_m_1_in), .ZN(n8) );
  LVT_XOR2HSV0 U5 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U6 ( .A1(n4), .A2(n7), .ZN(n5) );
endmodule


module cell_3_1947 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV1 U1 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_NAND2HSV1 U2 ( .A1(g_in), .A2(t_m_1_in), .ZN(n10) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_XOR2HSV0 U5 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_CLKNHSV0P5 U6 ( .I(n10), .ZN(n4) );
  LVT_NAND2HSV0P5 U7 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_INHSV0SR U8 ( .I(n9), .ZN(n5) );
endmodule


module cell_3_1946 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV1 U1 ( .A1(n4), .A2(n8), .B(n5), .ZN(t_i_out) );
  LVT_CLKNHSV2 U2 ( .I(n7), .ZN(n4) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U5 ( .A1(n8), .A2(n4), .ZN(n5) );
  LVT_NAND2HSV0 U6 ( .A1(g_in), .A2(t_m_1_in), .ZN(n8) );
endmodule


module cell_3_1945 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV1 U1 ( .A1(n4), .A2(n8), .B(n5), .ZN(t_i_out) );
  LVT_CLKNHSV0P5 U2 ( .I(n7), .ZN(n4) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U5 ( .A1(n8), .A2(n4), .ZN(n5) );
  LVT_NAND2HSV0 U6 ( .A1(g_in), .A2(t_m_1_in), .ZN(n8) );
endmodule


module cell_3_1944 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV0 U1 ( .A1(n4), .A2(n8), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(n8), .A2(n4), .ZN(n5) );
  LVT_INHSV2 U4 ( .I(n7), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0 U6 ( .A1(g_in), .A2(t_m_1_in), .ZN(n8) );
endmodule


module cell_3_1943 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n8), .B(n5), .ZN(t_i_out) );
  LVT_INHSV2 U2 ( .I(n7), .ZN(n4) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U5 ( .A1(n8), .A2(n4), .ZN(n5) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_1942 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n8), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(n8), .A2(n4), .ZN(n5) );
  LVT_INHSV2 U4 ( .I(n7), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0 U6 ( .A1(g_in), .A2(t_m_1_in), .ZN(n8) );
endmodule


module cell_3_1941 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_INAND2HSV2 U1 ( .A1(n9), .B1(n8), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n7), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U4 ( .A1(n9), .A2(n4), .ZN(n5) );
  LVT_NAND2HSV2 U5 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV0SR U6 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
endmodule


module cell_3_1940 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV0 U1 ( .A1(n4), .A2(n8), .B(n5), .ZN(t_i_out) );
  LVT_INHSV2 U2 ( .I(n7), .ZN(n4) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U5 ( .A1(n8), .A2(n4), .ZN(n5) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_1939 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV0 U1 ( .A1(n4), .A2(n8), .B(n5), .ZN(t_i_out) );
  LVT_INHSV2 U2 ( .I(n7), .ZN(n4) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U5 ( .A1(n8), .A2(n4), .ZN(n5) );
  LVT_NAND2HSV0 U6 ( .A1(g_in), .A2(t_m_1_in), .ZN(n8) );
endmodule


module cell_3_1938 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n8), .B(n5), .ZN(t_i_out) );
  LVT_INHSV2 U2 ( .I(n7), .ZN(n4) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U5 ( .A1(n8), .A2(n4), .ZN(n5) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_1937 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV0 U1 ( .A1(n4), .A2(n8), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(n8), .A2(n4), .ZN(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_INHSV2 U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(g_in), .A2(t_m_1_in), .ZN(n8) );
endmodule


module cell_3_1936 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_INAND2HSV2 U1 ( .A1(n9), .B1(n8), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n7), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U4 ( .A1(n9), .A2(n4), .ZN(n5) );
  LVT_CLKNAND2HSV0 U5 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV0SR U6 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
endmodule


module cell_3_1935 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_INAND2HSV2 U1 ( .A1(n9), .B1(n8), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n7), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U4 ( .A1(n9), .A2(n4), .ZN(n5) );
  LVT_CLKNAND2HSV0 U5 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV0SR U6 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
endmodule


module cell_3_1934 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV1 U1 ( .I(n10), .ZN(n4) );
  LVT_NAND2HSV2 U2 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_XOR2HSV0 U4 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_NAND2HSV0P5 U5 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0P5 U6 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_INHSV0SR U7 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV0 U8 ( .A1(g_in), .A2(t_m_1_in), .ZN(n10) );
endmodule


module cell_3_1933 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_INHSV2SR U2 ( .I(n8), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(g_in), .A2(t_m_1_in), .ZN(n8) );
  LVT_XOR2HSV0 U5 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U6 ( .A1(n4), .A2(n7), .ZN(n5) );
endmodule


module cell_3_1932 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_INHSV2SR U2 ( .I(n8), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(g_in), .A2(t_m_1_in), .ZN(n8) );
  LVT_XOR2HSV0 U5 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U6 ( .A1(n4), .A2(n7), .ZN(n5) );
endmodule


module cell_3_1931 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNHSV0 U1 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV0P5 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_INHSV1 U4 ( .I(n10), .ZN(n4) );
  LVT_NAND2HSV0 U5 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_XOR2HSV0 U6 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_NAND2HSV1 U7 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_NAND2HSV0 U8 ( .A1(g_in), .A2(t_m_1_in), .ZN(n10) );
endmodule


module cell_3_1930 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1929 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV1 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_INHSV2SR U2 ( .I(n8), .ZN(n4) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_1928 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_INHSV2 U2 ( .I(n8), .ZN(n4) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV0 U6 ( .A1(g_in), .A2(t_m_1_in), .ZN(n8) );
endmodule


module cell_3_1927 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(g_in), .A2(t_m_1_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1926 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1925 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1924 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module row_other_62 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_62 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_1954 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1953 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1952 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1951 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1950 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1949 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1948 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1947 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1946 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1945 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1944 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1943 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1942 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1941 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1940 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1939 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1938 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1937 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1936 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1935 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1934 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1933 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1932 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1931 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1930 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1929 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1928 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1927 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1926 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1925 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1924 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_2 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [31:0] a_in;
  input [31:0] g_in;
  input [31:0] b_in;
  input [31:0] t_m_1_in;
  input [30:0] t_i_1_in;
  input [30:0] t_i_2_in;
  output [31:0] a_out;
  output [31:0] g_out;
  output [30:0] t_i_1_out;
  output [30:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;
  wire   n1, n2, n4, n5, n7, n8, n10, n11, n13, n14, n16, n17, n19, n20, n22,
         n24, n26, n27;
  wire   [30:0] t0;
  wire   [30:0] t1;
  wire   [30:0] t2;
  wire   [30:0] t3;
  wire   [30:0] t4;
  wire   [30:0] t5;
  wire   [30:0] t6;
  wire   [30:0] t7;
  wire   [30:0] t8;
  wire   [30:0] t9;
  wire   [30:0] t10;
  wire   [30:0] t11;
  wire   [30:0] t12;
  wire   [30:0] t13;
  wire   [30:0] t14;
  wire   [30:0] t15;
  wire   [30:0] t16;
  wire   [30:0] t17;
  wire   [30:0] t18;
  wire   [30:0] t19;
  wire   [30:0] t20;
  wire   [30:0] t21;
  wire   [30:0] t22;
  wire   [30:0] t23;
  wire   [30:0] t24;
  wire   [30:0] t25;
  wire   [30:0] t26;
  wire   [30:0] t27;
  wire   [30:0] t28;
  wire   [30:0] t29;
  wire   [30:0] t30;
  assign a_out[30] = a_in[30];
  assign a_out[29] = a_in[29];
  assign a_out[28] = a_in[28];
  assign a_out[27] = a_in[27];
  assign a_out[26] = a_in[26];
  assign a_out[24] = a_in[24];
  assign a_out[21] = a_in[21];
  assign a_out[20] = a_in[20];
  assign a_out[19] = a_in[19];
  assign a_out[18] = a_in[18];
  assign a_out[17] = a_in[17];
  assign a_out[16] = a_in[16];
  assign a_out[15] = a_in[15];
  assign a_out[14] = a_in[14];
  assign a_out[13] = a_in[13];
  assign a_out[12] = a_in[12];
  assign a_out[11] = a_in[11];
  assign a_out[10] = a_in[10];
  assign a_out[9] = a_in[9];
  assign a_out[8] = a_in[8];
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[30] = g_in[30];
  assign g_out[29] = g_in[29];
  assign g_out[28] = g_in[28];
  assign g_out[27] = g_in[27];
  assign g_out[26] = g_in[26];
  assign g_out[21] = g_in[21];
  assign g_out[20] = g_in[20];
  assign g_out[19] = g_in[19];
  assign g_out[18] = g_in[18];
  assign g_out[17] = g_in[17];
  assign g_out[16] = g_in[16];
  assign g_out[15] = g_in[15];
  assign g_out[14] = g_in[14];
  assign g_out[13] = g_in[13];
  assign g_out[12] = g_in[12];
  assign g_out[11] = g_in[11];
  assign g_out[10] = g_in[10];
  assign g_out[9] = g_in[9];
  assign g_out[8] = g_in[8];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_2 u0 ( .a_in({a_in[31:26], n17, a_in[24], n8, n5, a_in[21:0]}), .g_in(
        {g_in[31:26], n20, n14, n11, n2, g_in[21:0]}), .b_in(b_in[31]), 
        .t_m_1_in(t_m_1_in[31]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(
        t_i_2_in), .t_i_1_out(t0), .t_i_2_out(t_i_2_out[30]) );
  row_other_92 u1 ( .a_in({a_in[31:26], a_out[25], a_in[24], a_out[23:22], 
        a_in[21:0]}), .g_in({g_in[31:26], g_out[25:22], g_in[21:0]}), .b_in(
        b_in[30]), .t_m_1_in(t_m_1_in[30]), .t_i_1_in(t0), .t_i_1_out(t1), 
        .t_i_2_out(t_i_2_out[29]) );
  row_other_91 u2 ( .a_in({a_in[31:26], a_out[25], a_in[24], a_out[23:22], 
        a_in[21:0]}), .g_in({g_in[31:26], g_out[25:22], g_in[21:0]}), .b_in(
        b_in[29]), .t_m_1_in(t_m_1_in[29]), .t_i_1_in(t1), .t_i_1_out(t2), 
        .t_i_2_out(t_i_2_out[28]) );
  row_other_90 u3 ( .a_in({a_in[31:26], a_out[25], a_in[24], a_out[23:22], 
        a_in[21:0]}), .g_in({g_in[31:26], g_out[25:22], g_in[21:0]}), .b_in(
        b_in[28]), .t_m_1_in(t_m_1_in[28]), .t_i_1_in(t2), .t_i_1_out(t3), 
        .t_i_2_out(t_i_2_out[27]) );
  row_other_89 u4 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[27]), .t_m_1_in(t_m_1_in[27]), 
        .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[26]) );
  row_other_88 u5 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[26]), .t_m_1_in(t_m_1_in[26]), 
        .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[25]) );
  row_other_87 u6 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[25]), .t_m_1_in(t_m_1_in[25]), 
        .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[24]) );
  row_other_86 u7 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[24]), .t_m_1_in(t_m_1_in[24]), 
        .t_i_1_in(t6), .t_i_1_out(t7), .t_i_2_out(t_i_2_out[23]) );
  row_other_85 u8 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[23]), .t_m_1_in(t_m_1_in[23]), 
        .t_i_1_in(t7), .t_i_1_out(t8), .t_i_2_out(t_i_2_out[22]) );
  row_other_84 u9 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[22]), .t_m_1_in(t_m_1_in[22]), 
        .t_i_1_in(t8), .t_i_1_out(t9), .t_i_2_out(t_i_2_out[21]) );
  row_other_83 u10 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[21]), .t_m_1_in(t_m_1_in[21]), 
        .t_i_1_in(t9), .t_i_1_out(t10), .t_i_2_out(t_i_2_out[20]) );
  row_other_82 u11 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[20]), .t_m_1_in(t_m_1_in[20]), 
        .t_i_1_in(t10), .t_i_1_out(t11), .t_i_2_out(t_i_2_out[19]) );
  row_other_81 u12 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[19]), .t_m_1_in(t_m_1_in[19]), 
        .t_i_1_in(t11), .t_i_1_out(t12), .t_i_2_out(t_i_2_out[18]) );
  row_other_80 u13 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[18]), .t_m_1_in(t_m_1_in[18]), 
        .t_i_1_in(t12), .t_i_1_out(t13), .t_i_2_out(t_i_2_out[17]) );
  row_other_79 u14 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[17]), .t_m_1_in(t_m_1_in[17]), 
        .t_i_1_in(t13), .t_i_1_out(t14), .t_i_2_out(t_i_2_out[16]) );
  row_other_78 u15 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[16]), .t_m_1_in(t_m_1_in[16]), 
        .t_i_1_in(t14), .t_i_1_out(t15), .t_i_2_out(t_i_2_out[15]) );
  row_other_77 u16 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[15]), .t_m_1_in(t_m_1_in[15]), 
        .t_i_1_in(t15), .t_i_1_out(t16), .t_i_2_out(t_i_2_out[14]) );
  row_other_76 u17 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[14]), .t_m_1_in(t_m_1_in[14]), 
        .t_i_1_in(t16), .t_i_1_out(t17), .t_i_2_out(t_i_2_out[13]) );
  row_other_75 u18 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[13]), .t_m_1_in(n27), 
        .t_i_1_in(t17), .t_i_1_out(t18), .t_i_2_out(t_i_2_out[12]) );
  row_other_74 u19 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[12]), .t_m_1_in(t_m_1_in[12]), 
        .t_i_1_in(t18), .t_i_1_out(t19), .t_i_2_out(t_i_2_out[11]) );
  row_other_73 u20 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[11]), .t_m_1_in(t_m_1_in[11]), 
        .t_i_1_in(t19), .t_i_1_out(t20), .t_i_2_out(t_i_2_out[10]) );
  row_other_72 u21 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[10]), .t_m_1_in(t_m_1_in[10]), 
        .t_i_1_in(t20), .t_i_1_out(t21), .t_i_2_out(t_i_2_out[9]) );
  row_other_71 u22 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[9]), .t_m_1_in(t_m_1_in[9]), 
        .t_i_1_in(t21), .t_i_1_out(t22), .t_i_2_out(t_i_2_out[8]) );
  row_other_70 u23 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[8]), .t_m_1_in(t_m_1_in[8]), 
        .t_i_1_in(t22), .t_i_1_out(t23), .t_i_2_out(t_i_2_out[7]) );
  row_other_69 u24 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[7]), .t_m_1_in(t_m_1_in[7]), 
        .t_i_1_in(t23), .t_i_1_out(t24), .t_i_2_out(t_i_2_out[6]) );
  row_other_68 u25 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[6]), .t_m_1_in(t_m_1_in[6]), 
        .t_i_1_in(t24), .t_i_1_out(t25), .t_i_2_out(t_i_2_out[5]) );
  row_other_67 u26 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[5]), .t_m_1_in(t_m_1_in[5]), 
        .t_i_1_in(t25), .t_i_1_out(t26), .t_i_2_out(t_i_2_out[4]) );
  row_other_66 u27 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[4]), .t_m_1_in(t_m_1_in[4]), 
        .t_i_1_in(t26), .t_i_1_out(t27), .t_i_2_out(t_i_2_out[3]) );
  row_other_65 u28 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[3]), .t_m_1_in(t_m_1_in[3]), 
        .t_i_1_in(t27), .t_i_1_out(t28), .t_i_2_out(t_i_2_out[2]) );
  row_other_64 u29 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[2]), .t_m_1_in(t_m_1_in[2]), 
        .t_i_1_in(t28), .t_i_1_out(t29), .t_i_2_out(t_i_2_out[1]) );
  row_other_63 u30 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[1]), .t_m_1_in(t_m_1_in[1]), 
        .t_i_1_in(t29), .t_i_1_out(t30), .t_i_2_out(t_i_2_out[0]) );
  row_other_62 u31 ( .a_in({a_out[31], a_in[30:26], a_out[25], a_in[24], 
        a_out[23:22], a_in[21:0]}), .g_in({g_out[31], g_in[30:26], 
        g_out[25:22], g_in[21:0]}), .b_in(b_in[0]), .t_m_1_in(t_m_1_in[0]), 
        .t_i_1_in(t30), .t_i_1_out(t_i_1_out), .t_i_2_out(t_i_1_out_0) );
  LVT_INHSV16SR U1 ( .I(n26), .ZN(n27) );
  LVT_CLKNHSV8 U2 ( .I(t_m_1_in[13]), .ZN(n26) );
  LVT_INHSV2 U3 ( .I(a_in[22]), .ZN(n4) );
  LVT_INHSV2 U4 ( .I(a_in[23]), .ZN(n7) );
  LVT_INHSV2 U5 ( .I(a_in[25]), .ZN(n16) );
  LVT_INHSV2 U6 ( .I(g_in[22]), .ZN(n1) );
  LVT_INHSV2 U7 ( .I(g_in[23]), .ZN(n10) );
  LVT_INHSV2 U8 ( .I(g_in[24]), .ZN(n13) );
  LVT_INHSV2 U9 ( .I(g_in[25]), .ZN(n19) );
  LVT_INHSV2SR U10 ( .I(n1), .ZN(n2) );
  LVT_INHSV2SR U11 ( .I(n1), .ZN(g_out[22]) );
  LVT_CLKNHSV2 U12 ( .I(n4), .ZN(n5) );
  LVT_INHSV2SR U13 ( .I(n4), .ZN(a_out[22]) );
  LVT_INHSV2 U14 ( .I(n7), .ZN(n8) );
  LVT_INHSV2SR U15 ( .I(n7), .ZN(a_out[23]) );
  LVT_CLKNHSV2 U16 ( .I(n10), .ZN(n11) );
  LVT_INHSV2SR U17 ( .I(n10), .ZN(g_out[23]) );
  LVT_CLKNHSV2 U18 ( .I(n13), .ZN(n14) );
  LVT_INHSV2SR U19 ( .I(n13), .ZN(g_out[24]) );
  LVT_INHSV2 U20 ( .I(n16), .ZN(n17) );
  LVT_INHSV2SR U21 ( .I(n16), .ZN(a_out[25]) );
  LVT_CLKNHSV2 U22 ( .I(n19), .ZN(n20) );
  LVT_INHSV2SR U23 ( .I(n19), .ZN(g_out[25]) );
  LVT_CLKNHSV4 U24 ( .I(n24), .ZN(g_out[31]) );
  LVT_INHSV0SR U25 ( .I(a_in[31]), .ZN(n22) );
  LVT_INHSV2 U26 ( .I(n22), .ZN(a_out[31]) );
  LVT_INHSV0SR U27 ( .I(g_in[31]), .ZN(n24) );
endmodule


module regist_32bit_13 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_32bit_12 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_31bit_8 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module PE_2 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro );
  input [31:0] a_in;
  input [31:0] g_in;
  input [31:0] b_in;
  input [30:0] t_i_1_in;
  input [30:0] t_i_2_in;
  output [31:0] a_out;
  output [31:0] g_out;
  output [31:0] b_out;
  output [30:0] t_i_1_out;
  output [30:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   n97, n98, n99, n100, l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] ,
         c_t_i_1_in_0, to_1, ti_1, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n40, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96;
  wire   [31:0] l_a;
  wire   [31:0] l_g;
  wire   [30:0] l_t_i_1_in;
  wire   [30:0] l_t_i_2_in;
  wire   [31:0] mux_b;
  wire   [31:0] mux_bq;
  wire   [30:0] to_7;
  wire   [30:0] ti_7;
  wire   [31:0] ao;
  wire   [31:0] go;
  wire   [30:0] to;

  LVT_AO22HSV0 U35 ( .A1(mux_bq[9]), .A2(n63), .B1(b_out[9]), .B2(n83), .Z(
        mux_b[9]) );
  LVT_AO22HSV0 U36 ( .A1(mux_bq[8]), .A2(n63), .B1(b_out[8]), .B2(n83), .Z(
        mux_b[8]) );
  LVT_AO22HSV0 U37 ( .A1(mux_bq[7]), .A2(n63), .B1(b_out[7]), .B2(n83), .Z(
        mux_b[7]) );
  LVT_AO22HSV0 U38 ( .A1(mux_bq[6]), .A2(n63), .B1(b_out[6]), .B2(n83), .Z(
        mux_b[6]) );
  LVT_AO22HSV0 U39 ( .A1(mux_bq[5]), .A2(n63), .B1(b_out[5]), .B2(n83), .Z(
        mux_b[5]) );
  LVT_AO22HSV0 U40 ( .A1(mux_bq[4]), .A2(n63), .B1(b_out[4]), .B2(n83), .Z(
        mux_b[4]) );
  LVT_AO22HSV0 U41 ( .A1(mux_bq[3]), .A2(n63), .B1(b_out[3]), .B2(n83), .Z(
        mux_b[3]) );
  LVT_AO22HSV0 U43 ( .A1(mux_bq[30]), .A2(n63), .B1(b_out[30]), .B2(n83), .Z(
        mux_b[30]) );
  LVT_AO22HSV0 U44 ( .A1(mux_bq[2]), .A2(n63), .B1(b_out[2]), .B2(n83), .Z(
        mux_b[2]) );
  LVT_AO22HSV0 U45 ( .A1(mux_bq[29]), .A2(n63), .B1(b_out[29]), .B2(n83), .Z(
        mux_b[29]) );
  LVT_AO22HSV0 U46 ( .A1(mux_bq[28]), .A2(n63), .B1(b_out[28]), .B2(n83), .Z(
        mux_b[28]) );
  LVT_AO22HSV0 U47 ( .A1(mux_bq[27]), .A2(n63), .B1(b_out[27]), .B2(n83), .Z(
        mux_b[27]) );
  LVT_AO22HSV0 U48 ( .A1(mux_bq[26]), .A2(n63), .B1(b_out[26]), .B2(n83), .Z(
        mux_b[26]) );
  LVT_AO22HSV0 U49 ( .A1(mux_bq[25]), .A2(n63), .B1(b_out[25]), .B2(n83), .Z(
        mux_b[25]) );
  LVT_AO22HSV0 U50 ( .A1(mux_bq[24]), .A2(n63), .B1(b_out[24]), .B2(n83), .Z(
        mux_b[24]) );
  LVT_AO22HSV0 U51 ( .A1(mux_bq[23]), .A2(n63), .B1(b_out[23]), .B2(n83), .Z(
        mux_b[23]) );
  LVT_AO22HSV0 U52 ( .A1(mux_bq[22]), .A2(n63), .B1(b_out[22]), .B2(n83), .Z(
        mux_b[22]) );
  LVT_AO22HSV0 U53 ( .A1(mux_bq[21]), .A2(n63), .B1(b_out[21]), .B2(n83), .Z(
        mux_b[21]) );
  LVT_AO22HSV0 U54 ( .A1(mux_bq[20]), .A2(n63), .B1(b_out[20]), .B2(n83), .Z(
        mux_b[20]) );
  LVT_AO22HSV0 U55 ( .A1(mux_bq[1]), .A2(n63), .B1(b_out[1]), .B2(n83), .Z(
        mux_b[1]) );
  LVT_AO22HSV0 U56 ( .A1(mux_bq[19]), .A2(n63), .B1(b_out[19]), .B2(n83), .Z(
        mux_b[19]) );
  LVT_AO22HSV0 U57 ( .A1(mux_bq[18]), .A2(n63), .B1(b_out[18]), .B2(n83), .Z(
        mux_b[18]) );
  LVT_AO22HSV0 U58 ( .A1(mux_bq[17]), .A2(n63), .B1(b_out[17]), .B2(n83), .Z(
        mux_b[17]) );
  LVT_AO22HSV0 U59 ( .A1(mux_bq[16]), .A2(n63), .B1(b_out[16]), .B2(n83), .Z(
        mux_b[16]) );
  LVT_AO22HSV0 U60 ( .A1(mux_bq[15]), .A2(n63), .B1(b_out[15]), .B2(n83), .Z(
        mux_b[15]) );
  LVT_AO22HSV0 U61 ( .A1(mux_bq[14]), .A2(n63), .B1(b_out[14]), .B2(n83), .Z(
        mux_b[14]) );
  LVT_AO22HSV0 U62 ( .A1(mux_bq[13]), .A2(n63), .B1(b_out[13]), .B2(n83), .Z(
        mux_b[13]) );
  LVT_AO22HSV0 U63 ( .A1(mux_bq[12]), .A2(n63), .B1(b_out[12]), .B2(n83), .Z(
        mux_b[12]) );
  LVT_AO22HSV0 U64 ( .A1(mux_bq[11]), .A2(n63), .B1(b_out[11]), .B2(n83), .Z(
        mux_b[11]) );
  LVT_AO22HSV0 U65 ( .A1(mux_bq[10]), .A2(n63), .B1(b_out[10]), .B2(n83), .Z(
        mux_b[10]) );
  LVT_AO22HSV0 U66 ( .A1(mux_bq[0]), .A2(n63), .B1(b_out[0]), .B2(n83), .Z(
        mux_b[0]) );
  LVT_NOR2HSV0 U67 ( .A1(n95), .A2(n83), .ZN(c_t_i_1_in_0) );
  LVT_AOI21HSV0 U69 ( .A1(n93), .A2(n92), .B(n83), .ZN(\c_t_i_1_in[0] ) );
  LVT_AND4HSV0 U71 ( .A1(n91), .A2(n90), .A3(n89), .A4(n88), .Z(n92) );
  LVT_NOR4HSV0 U72 ( .A1(l_t_i_1_in[9]), .A2(l_t_i_1_in[8]), .A3(l_t_i_1_in[7]), .A4(l_t_i_1_in[6]), .ZN(n88) );
  LVT_NOR4HSV0 U73 ( .A1(l_t_i_1_in[5]), .A2(l_t_i_1_in[4]), .A3(l_t_i_1_in[3]), .A4(l_t_i_1_in[30]), .ZN(n89) );
  LVT_NOR4HSV0 U74 ( .A1(l_t_i_1_in[2]), .A2(l_t_i_1_in[29]), .A3(
        l_t_i_1_in[28]), .A4(l_t_i_1_in[27]), .ZN(n90) );
  LVT_NOR4HSV0 U75 ( .A1(l_t_i_1_in[26]), .A2(l_t_i_1_in[25]), .A3(
        l_t_i_1_in[24]), .A4(l_t_i_1_in[23]), .ZN(n91) );
  LVT_AND4HSV0 U76 ( .A1(n87), .A2(n86), .A3(n85), .A4(n84), .Z(n93) );
  LVT_NOR4HSV0 U77 ( .A1(l_t_i_1_in[22]), .A2(l_t_i_1_in[21]), .A3(
        l_t_i_1_in[20]), .A4(l_t_i_1_in[1]), .ZN(n84) );
  LVT_NOR4HSV0 U78 ( .A1(l_t_i_1_in[19]), .A2(l_t_i_1_in[18]), .A3(
        l_t_i_1_in[17]), .A4(l_t_i_1_in[16]), .ZN(n85) );
  LVT_NOR4HSV0 U79 ( .A1(l_t_i_1_in[15]), .A2(l_t_i_1_in[14]), .A3(
        l_t_i_1_in[13]), .A4(l_t_i_1_in[12]), .ZN(n86) );
  LVT_NOR3HSV0 U80 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[11]), .A3(
        l_t_i_1_in[10]), .ZN(n87) );
  regist_32bit_17 u0 ( .clk(clk), .rstn(rstn), .in(a_in), .out(l_a) );
  regist_32bit_16 u1 ( .clk(clk), .rstn(rstn), .in(b_in), .out(b_out) );
  regist_32bit_15 u2 ( .clk(clk), .rstn(rstn), .in(g_in), .out(l_g) );
  regist_1bit_11 u3 ( .clk(clk), .rstn(rstn), .in(ctr), .out(l_ctr) );
  regist_1bit_10 u4 ( .clk(clk), .rstn(rstn), .in(n63), .out(ctro) );
  regist_31bit_11 u5 ( .clk(clk), .rstn(rstn), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_31bit_10 u6 ( .clk(clk), .rstn(rstn), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_9 u7 ( .clk(clk), .rstn(rstn), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_32bit_14 u9 ( .clk(clk), .rstn(rstn), .in(mux_b), .out(mux_bq) );
  regist_1bit_8 u10 ( .clk(clk), .rstn(rstn), .in(to_1), .out(ti_1) );
  regist_31bit_9 u11 ( .clk(clk), .rstn(rstn), .in({n75, n71, to_7[28:27], n44, 
        to_7[25:21], n61, to_7[19:13], n72, to_7[11:10], n26, to_7[8:3], n76, 
        n68, to_7[0]}), .out(ti_7) );
  PE_core_2 pe ( .a_in(l_a), .g_in(l_g), .b_in({n24, mux_bq[30:0]}), 
        .t_m_1_in({to_1, n75, n71, to_7[28:27], n44, to_7[25:21], n61, 
        to_7[19:13], n72, to_7[11:10], n26, to_7[8:3], n76, n68, to_7[0]}), 
        .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), 
        .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(
        go), .t_i_1_out(to), .t_i_2_out({t_i_2_out[30:27], n97, n98, 
        t_i_2_out[24:22], n99, t_i_2_out[20:10], n100, t_i_2_out[8:0]}), 
        .t_i_1_out_0(t_i_1_out_0) );
  regist_32bit_13 u12 ( .clk(clk), .rstn(rstn), .in(ao), .out(a_out) );
  regist_32bit_12 u13 ( .clk(clk), .rstn(rstn), .in(go), .out(g_out) );
  regist_31bit_8 u14 ( .clk(clk), .rstn(rstn), .in(to), .out(t_i_1_out) );
  LVT_INHSV5 U2 ( .I(n35), .ZN(n71) );
  LVT_NAND2HSV8 U3 ( .A1(n36), .A2(n37), .ZN(to_7[22]) );
  LVT_CLKNAND2HSV3 U4 ( .A1(t_i_2_out[7]), .A2(n96), .ZN(n18) );
  LVT_INHSV6 U5 ( .I(n30), .ZN(n75) );
  LVT_CLKNAND2HSV3 U6 ( .A1(n19), .A2(n20), .ZN(to_7[26]) );
  LVT_CLKNAND2HSV4 U7 ( .A1(n80), .A2(n79), .ZN(to_7[14]) );
  LVT_NAND2HSV4 U8 ( .A1(t_i_2_out[14]), .A2(n96), .ZN(n80) );
  LVT_OR2HSV12RD U9 ( .A1(n60), .A2(n59), .Z(to_7[15]) );
  LVT_NAND2HSV4 U10 ( .A1(t_i_2_out[8]), .A2(n96), .ZN(n58) );
  LVT_IAO22HSV4 U11 ( .B1(t_i_2_out[2]), .B2(n96), .A1(n34), .A2(n96), .ZN(n33) );
  LVT_CLKNAND2HSV2 U12 ( .A1(n97), .A2(n96), .ZN(n20) );
  LVT_AND2HSV4 U13 ( .A1(t_i_2_out[15]), .A2(n96), .Z(n60) );
  LVT_CLKNHSV10 U14 ( .I(n23), .ZN(n24) );
  LVT_INHSV4SR U15 ( .I(mux_bq[31]), .ZN(n23) );
  LVT_CLKNHSV8 U16 ( .I(n62), .ZN(n68) );
  LVT_NAND2HSV2 U17 ( .A1(ti_7[7]), .A2(ctro), .ZN(n17) );
  LVT_NAND2HSV2 U18 ( .A1(ti_7[10]), .A2(ctro), .ZN(n15) );
  LVT_CLKNAND2HSV4 U19 ( .A1(n54), .A2(n53), .ZN(to_7[4]) );
  LVT_NAND2HSV4 U20 ( .A1(n58), .A2(n57), .ZN(to_7[8]) );
  LVT_INHSV6 U21 ( .I(n43), .ZN(n44) );
  LVT_NAND2HSV2 U22 ( .A1(n56), .A2(n55), .ZN(to_7[6]) );
  LVT_INAND2HSV4 U23 ( .A1(n14), .B1(n22), .ZN(to_7[23]) );
  LVT_INHSV2 U24 ( .I(n21), .ZN(n14) );
  LVT_NAND2HSV8 U25 ( .A1(n70), .A2(n69), .ZN(to_7[28]) );
  LVT_IAO22HSV4 U26 ( .B1(t_i_2_out[20]), .B2(n96), .A1(n32), .A2(n96), .ZN(
        n31) );
  LVT_NAND2HSV4 U27 ( .A1(t_i_2_out[22]), .A2(n96), .ZN(n37) );
  LVT_OR2HSV12RD U28 ( .A1(n52), .A2(n51), .Z(to_7[17]) );
  LVT_CLKAND2HSV4 U29 ( .A1(t_i_2_out[0]), .A2(n96), .Z(n46) );
  LVT_INHSV3SR U30 ( .I(n31), .ZN(n61) );
  LVT_CLKNAND2HSV4 U31 ( .A1(t_i_2_out[10]), .A2(n96), .ZN(n16) );
  LVT_NAND2HSV4 U32 ( .A1(n15), .A2(n16), .ZN(to_7[10]) );
  LVT_INHSV12SR U33 ( .I(n25), .ZN(n26) );
  LVT_NAND2HSV4 U34 ( .A1(t_i_2_out[23]), .A2(n96), .ZN(n22) );
  LVT_NAND2HSV8 U42 ( .A1(n28), .A2(n27), .ZN(to_7[24]) );
  LVT_CLKNAND2HSV3 U68 ( .A1(t_i_2_out[24]), .A2(n96), .ZN(n28) );
  LVT_CLKNHSV6 U70 ( .I(l_ctr), .ZN(n94) );
  LVT_OR2HSV12RD U81 ( .A1(n46), .A2(n45), .Z(to_7[0]) );
  LVT_NAND2HSV4 U82 ( .A1(t_i_2_out[4]), .A2(n96), .ZN(n54) );
  LVT_CLKNHSV4 U83 ( .I(to_7[9]), .ZN(n25) );
  LVT_NAND2HSV3 U84 ( .A1(l_ctr), .A2(ti_1), .ZN(n81) );
  LVT_CLKNAND2HSV8 U85 ( .A1(n94), .A2(l_t_i_1_in_0), .ZN(n82) );
  LVT_CLKNAND2HSV8 U86 ( .A1(n81), .A2(n82), .ZN(to_1) );
  LVT_INHSV4SR U87 ( .I(to_7[26]), .ZN(n43) );
  LVT_NAND2HSV4 U88 ( .A1(n17), .A2(n18), .ZN(to_7[7]) );
  LVT_CLKAND2HSV4 U89 ( .A1(t_i_2_out[11]), .A2(n96), .Z(n50) );
  LVT_CLKNAND2HSV3 U90 ( .A1(t_i_2_out[27]), .A2(n96), .ZN(n65) );
  LVT_NAND2HSV4 U91 ( .A1(n64), .A2(n65), .ZN(to_7[27]) );
  LVT_OR2HSV16RD U92 ( .A1(n48), .A2(n47), .Z(to_7[21]) );
  LVT_AND2HSV8 U93 ( .A1(n99), .A2(n96), .Z(n48) );
  LVT_INHSV4SR U94 ( .I(n33), .ZN(n76) );
  LVT_NAND2HSV2 U95 ( .A1(t_i_2_out[6]), .A2(n96), .ZN(n56) );
  LVT_INHSV2 U96 ( .I(ti_7[2]), .ZN(n34) );
  LVT_OR2HSV12RD U97 ( .A1(n67), .A2(n66), .Z(to_7[5]) );
  LVT_CLKAND2HSV4 U98 ( .A1(t_i_2_out[5]), .A2(n96), .Z(n67) );
  LVT_INHSV6 U99 ( .I(ctro), .ZN(n96) );
  LVT_INHSV2 U100 ( .I(n29), .ZN(n83) );
  LVT_INHSV2 U101 ( .I(ti_7[20]), .ZN(n32) );
  LVT_NAND2HSV2 U102 ( .A1(ti_7[26]), .A2(ctro), .ZN(n19) );
  LVT_NAND2HSV2 U103 ( .A1(ti_7[23]), .A2(ctro), .ZN(n21) );
  LVT_NAND2HSV2 U104 ( .A1(ti_7[24]), .A2(ctro), .ZN(n27) );
  LVT_OR2HSV12RD U105 ( .A1(n50), .A2(n49), .Z(to_7[11]) );
  LVT_INHSV2 U106 ( .I(n83), .ZN(n63) );
  LVT_INHSV0SR U107 ( .I(n94), .ZN(n29) );
  LVT_AOI22HSV4 U108 ( .A1(ti_7[30]), .A2(ctro), .B1(t_i_2_out[30]), .B2(n96), 
        .ZN(n30) );
  LVT_INHSV4SR U109 ( .I(n42), .ZN(n72) );
  LVT_CLKNAND2HSV3 U110 ( .A1(t_i_2_out[28]), .A2(n96), .ZN(n70) );
  LVT_AOI22HSV4 U111 ( .A1(ti_7[29]), .A2(ctro), .B1(t_i_2_out[29]), .B2(n96), 
        .ZN(n35) );
  LVT_NAND2HSV2 U112 ( .A1(ti_7[22]), .A2(ctro), .ZN(n36) );
  LVT_INHSV0SR U113 ( .I(n99), .ZN(n38) );
  LVT_INHSV2 U114 ( .I(n38), .ZN(t_i_2_out[21]) );
  LVT_INHSV0SR U115 ( .I(n98), .ZN(n40) );
  LVT_INHSV2 U116 ( .I(n40), .ZN(t_i_2_out[25]) );
  LVT_AOI22HSV4 U117 ( .A1(ti_7[12]), .A2(ctro), .B1(t_i_2_out[12]), .B2(n96), 
        .ZN(n42) );
  LVT_AND2HSV0RD U118 ( .A1(ti_7[0]), .A2(ctro), .Z(n45) );
  LVT_AND2HSV0RD U119 ( .A1(ti_7[21]), .A2(ctro), .Z(n47) );
  LVT_AND2HSV0RD U120 ( .A1(ti_7[11]), .A2(ctro), .Z(n49) );
  LVT_AND2HSV0RD U121 ( .A1(ti_7[17]), .A2(ctro), .Z(n51) );
  LVT_AND2HSV8 U122 ( .A1(t_i_2_out[17]), .A2(n96), .Z(n52) );
  LVT_NAND2HSV0P5 U123 ( .A1(ti_7[4]), .A2(ctro), .ZN(n53) );
  LVT_NAND2HSV0 U124 ( .A1(ti_7[6]), .A2(ctro), .ZN(n55) );
  LVT_NAND2HSV0 U125 ( .A1(ti_7[8]), .A2(ctro), .ZN(n57) );
  LVT_AND2HSV0RD U126 ( .A1(ti_7[15]), .A2(ctro), .Z(n59) );
  LVT_AOI22HSV4 U127 ( .A1(ti_7[1]), .A2(ctro), .B1(t_i_2_out[1]), .B2(n96), 
        .ZN(n62) );
  LVT_AO22HSV1 U128 ( .A1(n24), .A2(n63), .B1(b_out[31]), .B2(n83), .Z(
        mux_b[31]) );
  LVT_NAND2HSV0 U129 ( .A1(ti_7[27]), .A2(ctro), .ZN(n64) );
  LVT_AND2HSV0RD U130 ( .A1(ti_7[5]), .A2(ctro), .Z(n66) );
  LVT_NAND2HSV0 U131 ( .A1(ti_7[28]), .A2(ctro), .ZN(n69) );
  LVT_INHSV0SR U132 ( .I(n100), .ZN(n73) );
  LVT_INHSV2 U133 ( .I(n73), .ZN(t_i_2_out[9]) );
  LVT_AO22HSV4 U134 ( .A1(ti_7[16]), .A2(ctro), .B1(t_i_2_out[16]), .B2(n96), 
        .Z(to_7[16]) );
  LVT_AO22HSV4 U135 ( .A1(ti_7[18]), .A2(ctro), .B1(t_i_2_out[18]), .B2(n96), 
        .Z(to_7[18]) );
  LVT_AO22HSV4 U136 ( .A1(ti_7[13]), .A2(ctro), .B1(t_i_2_out[13]), .B2(n96), 
        .Z(to_7[13]) );
  LVT_INHSV0SR U137 ( .I(n97), .ZN(n77) );
  LVT_INHSV2 U138 ( .I(n77), .ZN(t_i_2_out[26]) );
  LVT_NAND2HSV0 U139 ( .A1(ti_7[14]), .A2(ctro), .ZN(n79) );
  LVT_AO22HSV4 U140 ( .A1(ti_7[19]), .A2(ctro), .B1(t_i_2_out[19]), .B2(n96), 
        .Z(to_7[19]) );
  LVT_AO22HSV4 U141 ( .A1(ti_7[3]), .A2(ctro), .B1(t_i_2_out[3]), .B2(n96), 
        .Z(to_7[3]) );
  LVT_AO22HSV4 U142 ( .A1(ti_7[25]), .A2(ctro), .B1(n98), .B2(n96), .Z(
        to_7[25]) );
  LVT_AO22HSV4 U143 ( .A1(ti_7[9]), .A2(ctro), .B1(n100), .B2(n96), .Z(to_7[9]) );
  LVT_INHSV1 U144 ( .I(l_t_i_1_in_0), .ZN(n95) );
endmodule


module regist_32bit_11 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV4 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV4 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV4 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV4 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV4 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV4 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV4 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV4 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV4 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n2), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n2), .Q(out[31]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n1), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n1), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n1), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n1), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n1), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n1), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n1), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n2), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n2), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n2), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_CLKNHSV4 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_32bit_10 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV2 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n2), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n2), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n2), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_32bit_9 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV4 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n2), .Q(out[31]) );
  LVT_DRNQHSV4 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV4 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV4 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV4 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV4 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV4 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n2), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n1), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n1), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n1), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n1), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n1), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n1), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n1), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n2), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n2), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n2), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_CLKNHSV4 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_1bit_7 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_6 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_31bit_7 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n1), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n1), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n1), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n1), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n1), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n1), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n1), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n2) );
  LVT_CLKNHSV4 U4 ( .I(n2), .ZN(n1) );
endmodule


module regist_31bit_6 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n1), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(rstn), .Q(out[27])
         );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n1), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n1), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(rstn), .Q(out[28])
         );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n1), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n1), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n1), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n1), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n2) );
  LVT_CLKNHSV4 U4 ( .I(n2), .ZN(n1) );
endmodule


module regist_1bit_5 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_32bit_8 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV4 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n2), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n2), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n2), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n2), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n2), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n2), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n2), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_CLKNHSV4 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_1bit_4 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_31bit_5 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n2), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n2), .Q(out[28]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n2), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n2), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n2), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n2), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n1) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n2) );
endmodule


module cell_3_1923 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_61 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_60 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_59 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_58 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_57 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_56 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_55 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_54 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_53 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_52 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_51 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_50 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_49 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_48 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_47 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_46 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_45 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_44 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_43 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_42 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_41 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_NAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_4_40 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_39 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_38 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_37 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_36 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_35 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_34 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_33 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV2 U1 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_32 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
endmodule


module cell_4_31 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12;

  LVT_INHSV3SR U1 ( .I(n10), .ZN(n2) );
  LVT_IOA21HSV4 U2 ( .A1(n9), .A2(n10), .B(n3), .ZN(t_i_out) );
  LVT_CLKNHSV2 U3 ( .I(n12), .ZN(n6) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n2), .A2(n1), .ZN(n3) );
  LVT_NAND2HSV0 U5 ( .A1(n11), .A2(n12), .ZN(n7) );
  LVT_CLKNAND2HSV3 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n12) );
  LVT_NAND2HSV2 U7 ( .A1(n7), .A2(n8), .ZN(n10) );
  LVT_CLKNHSV0P5 U8 ( .I(n11), .ZN(n5) );
  LVT_NAND2HSV2 U9 ( .A1(n5), .A2(n6), .ZN(n8) );
  LVT_CLKAND2HSV1 U10 ( .A1(b_in), .A2(a_in), .Z(n11) );
  LVT_INHSV2 U11 ( .I(n9), .ZN(n1) );
  LVT_XNOR2HSV1 U12 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n9) );
endmodule


module row_1_1 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [31:0] t_i_1_in;
  input [30:0] t_i_2_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_3_1923 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_61 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(t_i_1_out[1])
         );
  cell_4_60 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(t_i_1_out[2])
         );
  cell_4_59 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(t_i_1_out[3])
         );
  cell_4_58 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(t_i_1_out[4])
         );
  cell_4_57 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(t_i_1_out[5])
         );
  cell_4_56 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(t_i_1_out[6])
         );
  cell_4_55 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(t_i_1_out[7])
         );
  cell_4_54 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_2_in(t_i_2_in[7]), .t_i_out(t_i_1_out[8])
         );
  cell_4_53 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[9]), .t_i_2_in(t_i_2_in[8]), .t_i_out(t_i_1_out[9])
         );
  cell_4_52 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[10]), .t_i_2_in(t_i_2_in[9]), .t_i_out(
        t_i_1_out[10]) );
  cell_4_51 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[11]), .t_i_2_in(t_i_2_in[10]), .t_i_out(
        t_i_1_out[11]) );
  cell_4_50 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[12]), .t_i_2_in(t_i_2_in[11]), .t_i_out(
        t_i_1_out[12]) );
  cell_4_49 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[13]), .t_i_2_in(t_i_2_in[12]), .t_i_out(
        t_i_1_out[13]) );
  cell_4_48 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[14]), .t_i_2_in(t_i_2_in[13]), .t_i_out(
        t_i_1_out[14]) );
  cell_4_47 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[15]), .t_i_2_in(t_i_2_in[14]), .t_i_out(
        t_i_1_out[15]) );
  cell_4_46 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[16]), .t_i_2_in(t_i_2_in[15]), .t_i_out(
        t_i_1_out[16]) );
  cell_4_45 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[17]), .t_i_2_in(t_i_2_in[16]), .t_i_out(
        t_i_1_out[17]) );
  cell_4_44 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[18]), .t_i_2_in(t_i_2_in[17]), .t_i_out(
        t_i_1_out[18]) );
  cell_4_43 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[19]), .t_i_2_in(t_i_2_in[18]), .t_i_out(
        t_i_1_out[19]) );
  cell_4_42 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[20]), .t_i_2_in(t_i_2_in[19]), .t_i_out(
        t_i_1_out[20]) );
  cell_4_41 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_2_in(t_i_2_in[20]), .t_i_out(
        t_i_1_out[21]) );
  cell_4_40 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_2_in(t_i_2_in[21]), .t_i_out(
        t_i_1_out[22]) );
  cell_4_39 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_2_in(t_i_2_in[22]), .t_i_out(
        t_i_1_out[23]) );
  cell_4_38 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_2_in(t_i_2_in[23]), .t_i_out(
        t_i_1_out[24]) );
  cell_4_37 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_2_in(t_i_2_in[24]), .t_i_out(
        t_i_1_out[25]) );
  cell_4_36 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_2_in(t_i_2_in[25]), .t_i_out(
        t_i_1_out[26]) );
  cell_4_35 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_2_in(t_i_2_in[26]), .t_i_out(
        t_i_1_out[27]) );
  cell_4_34 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_2_in(t_i_2_in[27]), .t_i_out(
        t_i_1_out[28]) );
  cell_4_33 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_2_in(t_i_2_in[28]), .t_i_out(
        t_i_1_out[29]) );
  cell_4_32 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_2_in(t_i_2_in[29]), .t_i_out(
        t_i_1_out[30]) );
  cell_4_31 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[31]), .t_i_2_in(t_i_2_in[30]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV2 U1 ( .I(n2), .ZN(n3) );
  LVT_INHSV2 U2 ( .I(n2), .ZN(n1) );
  LVT_INHSV0SR U3 ( .I(t_m_1_in), .ZN(n2) );
endmodule


module cell_2_61 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1922 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1921 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1920 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1919 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1918 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1917 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1916 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1915 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1914 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1913 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1912 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1911 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1910 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1909 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1908 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1907 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1906 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1905 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1904 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1903 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1902 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1901 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1900 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1899 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1898 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1897 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_1896 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1895 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1894 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1893 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_1892 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12;

  LVT_NAND2HSV0P5 U1 ( .A1(n12), .A2(n10), .ZN(n5) );
  LVT_CLKNHSV2 U2 ( .I(n12), .ZN(n2) );
  LVT_CLKNAND2HSV3 U3 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n12) );
  LVT_NAND2HSV2 U5 ( .A1(n8), .A2(n9), .ZN(n10) );
  LVT_INAND2HSV2 U6 ( .A1(n11), .B1(n7), .ZN(n9) );
  LVT_NAND2HSV2 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2SR U8 ( .I(n10), .ZN(n4) );
  LVT_INHSV2 U9 ( .I(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV0P5 U10 ( .A1(t_i_1_in), .A2(n11), .ZN(n8) );
  LVT_NAND2HSV0 U11 ( .A1(b_in), .A2(a_in), .ZN(n11) );
endmodule


module row_other_61 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_61 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1922 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1921 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1920 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1919 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1918 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1917 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1916 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1915 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1914 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1913 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1912 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1911 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1910 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1909 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1908 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1907 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1906 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1905 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1904 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1903 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1902 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1901 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1900 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1899 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1898 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1897 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1896 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1895 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1894 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1893 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1892 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV3SR U1 ( .I(n2), .ZN(n1) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n2) );
  LVT_BUFHSV2RT U3 ( .I(n1), .Z(n3) );
endmodule


module cell_2_60 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1891 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1890 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1889 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1888 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1887 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1886 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1885 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1884 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1883 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1882 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1881 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1880 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1879 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1878 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1877 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1876 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1875 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1874 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1873 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1872 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1871 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1870 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1869 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1868 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1867 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1866 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1865 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1864 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1863 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1862 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1861 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV4 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNHSV2 U2 ( .I(n9), .ZN(n2) );
  LVT_INHSV4 U4 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV4 U5 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV2 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV4 U7 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV0P5 U8 ( .A1(n9), .A2(n7), .ZN(n5) );
endmodule


module row_other_60 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_60 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1891 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1890 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1889 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1888 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1887 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1886 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1885 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1884 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1883 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1882 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1881 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1880 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1879 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1878 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1877 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1876 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1875 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1874 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1873 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1872 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1871 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1870 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1869 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1868 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1867 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1866 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1865 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1864 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1863 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1862 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1861 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV4 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_59 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_1860 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1859 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1858 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1857 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1856 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1855 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1854 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1853 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1852 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1851 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1850 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1849 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1848 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1847 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1846 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1845 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1844 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1843 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1842 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1841 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1840 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1839 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1838 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1837 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1836 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1835 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1834 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1833 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0P5 U4 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_CLKNHSV0P5 U5 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_1832 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1831 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_INHSV2P5 U1 ( .I(n8), .ZN(n4) );
  LVT_CLKNAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U4 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV2 U5 ( .A1(n7), .A2(n4), .ZN(n5) );
  LVT_XOR2HSV4 U6 ( .A1(t_i_1_in), .A2(n6), .Z(n7) );
endmodule


module cell_3_1830 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4, n5, n6, n7, n8;

  LVT_INHSV3SR U1 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV4 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XNOR2HSV4 U3 ( .A1(t_i_1_in), .A2(n2), .ZN(n3) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV4 U5 ( .A1(n4), .A2(n3), .ZN(n6) );
  LVT_XOR2HSV0 U6 ( .A1(t_i_1_in), .A2(n2), .Z(n7) );
  LVT_CLKNAND2HSV1 U7 ( .A1(n8), .A2(n7), .ZN(n5) );
  LVT_CLKAND2HSV2 U8 ( .A1(b_in), .A2(a_in), .Z(n2) );
endmodule


module row_other_59 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_59 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1860 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1859 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1858 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1857 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1856 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1855 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1854 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1853 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1852 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1851 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1850 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1849 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1848 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1847 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1846 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1845 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1844 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1843 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1842 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1841 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1840 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1839 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1838 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1837 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1836 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1835 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1834 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1833 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1832 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1831 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1830 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV2 U1 ( .I(t_m_1_in), .ZN(n2) );
  LVT_CLKNHSV4 U2 ( .I(n2), .ZN(n1) );
  LVT_INHSV0SR U3 ( .I(n2), .ZN(n3) );
endmodule


module cell_2_58 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1829 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1828 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1827 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1826 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1825 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1824 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1823 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1822 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1821 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1820 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1819 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1818 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1817 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1816 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1815 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1814 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1813 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1812 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1811 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1810 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1809 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1808 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1807 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1806 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1805 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1804 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1803 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1802 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1801 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_1800 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV3 U1 ( .A1(n4), .A2(n2), .ZN(n6) );
  LVT_NAND2HSV2 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_XOR2HSV0 U3 ( .A1(n8), .A2(t_i_1_in), .Z(n2) );
  LVT_NAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV0P5 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2 U7 ( .I(n9), .ZN(n4) );
  LVT_XNOR2HSV1 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module cell_3_1799 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_58 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_58 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1829 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1828 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1827 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1826 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1825 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1824 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1823 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1822 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1821 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1820 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1819 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1818 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1817 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1816 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1815 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1814 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1813 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1812 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1811 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1810 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1809 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1808 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1807 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1806 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1805 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1804 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1803 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1802 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1801 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1800 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1799 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV4 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_57 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1798 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1797 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1796 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1795 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1794 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1793 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1792 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1791 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1790 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1789 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1788 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1787 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1786 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1785 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1784 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1783 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1782 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1781 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1780 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1779 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1778 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1777 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1776 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1775 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1774 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1773 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1772 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1771 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1770 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1769 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_1768 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_INHSV3SR U4 ( .I(n9), .ZN(n5) );
  LVT_CLKNAND2HSV3 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_CLKXOR2HSV4 U6 ( .A1(t_i_1_in), .A2(n8), .Z(n9) );
  LVT_INHSV2 U7 ( .I(n10), .ZN(n4) );
  LVT_NAND2HSV2 U8 ( .A1(n4), .A2(n9), .ZN(n7) );
endmodule


module row_other_57 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4, n5;

  cell_2_57 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1798 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1797 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1796 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1795 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1794 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1793 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1792 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1791 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n5), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1790 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1789 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1788 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1787 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1786 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1785 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1784 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1783 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1782 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1781 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1780 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1779 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1778 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1777 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1776 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1775 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1774 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1773 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1772 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1771 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1770 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1769 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1768 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV2 U1 ( .I(n1), .ZN(n3) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
  LVT_INHSV0SR U3 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(n4), .ZN(n5) );
  LVT_INHSV0SR U5 ( .I(n3), .ZN(n4) );
endmodule


module cell_2_56 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1767 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1766 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1765 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1764 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1763 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1762 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1761 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1760 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1759 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1758 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1757 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1756 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1755 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1754 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1753 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1752 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1751 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1750 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1749 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1748 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1747 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1746 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1745 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1744 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1743 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1742 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1741 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U3 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV0 U5 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_3_1740 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1739 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1738 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_1737 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2SR U4 ( .I(n9), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV2 U6 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U7 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
  LVT_NAND2HSV0P5 U8 ( .A1(n9), .A2(n7), .ZN(n5) );
endmodule


module row_other_56 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_56 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1767 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1766 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1765 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1764 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1763 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1762 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1761 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1760 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1759 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1758 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1757 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1756 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1755 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1754 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1753 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1752 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1751 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1750 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1749 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1748 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1747 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1746 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1745 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1744 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1743 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1742 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1741 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1740 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1739 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1738 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1737 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKBUFHSV4 U1 ( .I(t_m_1_in), .Z(n2) );
  LVT_BUFHSV8 U2 ( .I(n2), .Z(n1) );
endmodule


module cell_2_55 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1736 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1735 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1734 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1733 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1732 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1731 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1730 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1729 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1728 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1727 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1726 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1725 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1724 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1723 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1722 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1721 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1720 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1719 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1718 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1717 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1716 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1715 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1714 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1713 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1712 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1711 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1710 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1709 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1708 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1707 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_1706 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n7), .A2(n5), .ZN(n4) );
  LVT_CLKNAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n7) );
  LVT_OAI21HSV2 U4 ( .A1(n2), .A2(n5), .B(n4), .ZN(t_i_out) );
  LVT_NAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_XNOR2HSV4 U6 ( .A1(t_i_1_in), .A2(n6), .ZN(n5) );
endmodule


module row_other_55 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_55 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_1736 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1735 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1734 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1733 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1732 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1731 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1730 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1729 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1728 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1727 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1726 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1725 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1724 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1723 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1722 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1721 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1720 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1719 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1718 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1717 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1716 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1715 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1714 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1713 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1712 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1711 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1710 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1709 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1708 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1707 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1706 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_54 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_1705 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1704 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1703 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1702 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1701 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1700 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1699 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1698 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1697 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1696 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1695 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1694 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1693 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1692 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1691 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1690 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1689 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1688 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1687 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1686 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1685 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1684 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1683 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1682 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1681 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1680 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1679 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1678 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INAND2HSV2 U2 ( .A1(n9), .B1(n8), .ZN(n6) );
  LVT_NAND2HSV0P5 U4 ( .A1(n9), .A2(n4), .ZN(n5) );
  LVT_NAND2HSV2 U5 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNHSV2 U6 ( .I(n8), .ZN(n4) );
  LVT_XOR2HSV2 U7 ( .A1(n7), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_3_1677 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1676 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_CLKXOR2HSV2 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_1675 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV2 U5 ( .I(n7), .ZN(n4) );
  LVT_INHSV2 U6 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV2 U7 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_54 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_2_54 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1705 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1704 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1703 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1702 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1701 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1700 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1699 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1698 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1697 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1696 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1695 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1694 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1693 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1692 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1691 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1690 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1689 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1688 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1687 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1686 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1685 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1684 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1683 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1682 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1681 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1680 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1679 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1678 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1677 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1676 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1675 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV20 U1 ( .I(n1), .ZN(n2) );
  LVT_CLKNHSV8 U2 ( .I(n4), .ZN(n1) );
  LVT_INHSV3SR U3 ( .I(n3), .ZN(n4) );
  LVT_INHSV0SR U4 ( .I(t_m_1_in), .ZN(n3) );
endmodule


module cell_2_53 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1674 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1673 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1672 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1671 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1670 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1669 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1668 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1667 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1666 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1665 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1664 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1663 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1662 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1661 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1660 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1659 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1658 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1657 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1656 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1655 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1654 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1653 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1652 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1651 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1650 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1649 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1648 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1647 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1646 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1645 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1644 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_53 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1;

  cell_2_53 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1674 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1673 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1672 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1671 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1670 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1669 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1668 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1667 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1666 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1665 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1664 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1663 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1662 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1661 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1660 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1659 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1658 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1657 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1656 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1655 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1654 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1653 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1652 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1651 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1650 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1649 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1648 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1647 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1646 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1645 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1644 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV16RT U1 ( .I(t_m_1_in), .Z(n1) );
endmodule


module cell_2_52 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1643 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1642 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1641 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1640 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1639 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1638 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1637 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1636 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1635 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1634 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1633 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1632 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1631 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1630 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1629 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1628 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1627 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1626 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1625 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1624 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1623 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1622 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1621 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1620 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1619 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1618 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1617 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1616 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1615 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1614 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1613 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_52 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_52 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1643 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1642 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1641 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1640 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1639 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1638 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1637 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1636 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1635 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1634 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1633 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1632 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1631 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1630 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1629 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1628 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1627 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1626 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1625 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1624 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1623 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1622 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1621 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1620 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1619 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1618 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1617 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1616 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1615 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1614 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1613 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV4RT U1 ( .I(t_m_1_in), .Z(n1) );
  LVT_INHSV6SR U2 ( .I(n2), .ZN(n3) );
  LVT_CLKNHSV2 U3 ( .I(t_m_1_in), .ZN(n2) );
endmodule


module cell_2_51 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1612 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1611 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1610 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1609 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1608 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1607 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1606 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1605 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1604 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1603 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1602 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1601 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1600 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1599 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1598 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1597 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1596 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1595 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1594 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1593 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1592 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1591 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1590 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1589 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1588 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1587 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1586 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1585 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1584 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1583 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_CLKNHSV2 U5 ( .I(n10), .ZN(n4) );
  LVT_INHSV0SR U6 ( .I(n9), .ZN(n5) );
  LVT_XOR2HSV2 U7 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_NAND2HSV0P5 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_1582 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_51 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1;

  cell_2_51 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1612 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1611 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1610 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1609 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1608 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1607 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1606 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1605 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1604 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1603 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1602 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1601 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1600 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1599 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1598 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1597 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1596 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1595 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1594 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1593 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1592 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1591 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1590 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1589 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1588 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1587 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1586 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1585 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1584 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1583 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1582 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV2 U1 ( .I(t_m_1_in), .Z(n1) );
endmodule


module cell_2_50 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1581 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1580 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1579 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1578 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1577 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1576 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1575 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1574 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1573 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1572 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1571 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1570 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1569 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1568 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1567 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1566 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1565 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1564 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1563 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1562 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1561 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1560 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1559 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1558 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1557 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1556 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1555 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1554 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1553 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1552 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1551 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV2 U1 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_CLKNAND2HSV1 U2 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_NAND2HSV4 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_CLKNHSV0 U6 ( .I(n9), .ZN(n5) );
  LVT_INHSV3SR U7 ( .I(n10), .ZN(n4) );
  LVT_NAND2HSV0P5 U8 ( .A1(n10), .A2(n5), .ZN(n6) );
endmodule


module row_other_50 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_2_50 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1581 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1580 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1579 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1578 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1577 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1576 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1575 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1574 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1573 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1572 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1571 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1570 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1569 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1568 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1567 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1566 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1565 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1564 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1563 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1562 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1561 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1560 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1559 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1558 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1557 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1556 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1555 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1554 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1553 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1552 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1551 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV5 U1 ( .I(n3), .ZN(n4) );
  LVT_INHSV2 U2 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U3 ( .I(n4), .ZN(n2) );
  LVT_CLKNHSV0P5 U4 ( .I(t_m_1_in), .ZN(n3) );
endmodule


module cell_2_49 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1550 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1549 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1548 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1547 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1546 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1545 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1544 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1543 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1542 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1541 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1540 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1539 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1538 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1537 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1536 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1535 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1534 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1533 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1532 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1531 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1530 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1529 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1528 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1527 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1526 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1525 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U5 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0P5 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_1524 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1523 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1522 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1521 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1520 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_49 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_49 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1550 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1549 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1548 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1547 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1546 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1545 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1544 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1543 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1542 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1541 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1540 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1539 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1538 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1537 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1536 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1535 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1534 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1533 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1532 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1531 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1530 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1529 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1528 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1527 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1526 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1525 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1524 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1523 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1522 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1521 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1520 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV6 U1 ( .I(n2), .ZN(n3) );
  LVT_INHSV6 U2 ( .I(t_m_1_in), .ZN(n2) );
  LVT_BUFHSV2RT U3 ( .I(n3), .Z(n1) );
endmodule


module cell_2_48 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1519 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1518 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1517 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1516 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1515 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1514 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1513 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1512 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1511 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1510 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1509 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1508 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1507 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1506 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1505 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1504 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1503 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1502 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_1501 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1500 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1499 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1498 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1497 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1496 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1495 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1494 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1493 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1492 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1491 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1490 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_INHSV2SR U1 ( .I(n8), .ZN(n4) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV0P5 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XOR2HSV2 U6 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
endmodule


module cell_3_1489 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_48 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1;

  cell_2_48 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1519 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1518 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1517 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1516 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1515 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1514 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1513 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1512 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1511 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1510 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1509 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1508 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1507 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1506 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1505 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1504 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1503 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1502 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1501 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1500 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1499 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1498 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1497 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1496 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1495 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1494 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1493 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1492 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1491 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1490 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1489 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV2 U1 ( .I(t_m_1_in), .Z(n1) );
endmodule


module cell_2_47 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1488 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1487 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1486 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1485 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1484 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1483 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1482 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1481 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1480 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1479 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1478 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1477 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1476 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1475 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1474 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1473 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1472 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1471 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1470 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1469 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1468 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1467 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1466 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1465 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1464 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1463 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1462 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1461 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1460 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1459 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1458 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n2), .A2(n4), .ZN(n5) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNHSV2P5 U4 ( .I(n9), .ZN(n2) );
  LVT_CLKNHSV2P5 U5 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV2 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV0P5 U7 ( .A1(n9), .A2(n7), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_47 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_2_47 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1488 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1487 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1486 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1485 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1484 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1483 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1482 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1481 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1480 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1479 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1478 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1477 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1476 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1475 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1474 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1473 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1472 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1471 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1470 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1469 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1468 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1467 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1466 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1465 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1464 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1463 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1462 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1461 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1460 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1459 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1458 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV2 U1 ( .I(t_m_1_in), .ZN(n3) );
  LVT_INHSV6 U2 ( .I(n3), .ZN(n4) );
  LVT_INHSV0SR U3 ( .I(n4), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_46 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_1457 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1456 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1455 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1454 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1453 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1452 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1451 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1450 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1449 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1448 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1447 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1446 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1445 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1444 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1443 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1442 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1441 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1440 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1439 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1438 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1437 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1436 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1435 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1434 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1433 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1432 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1431 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1430 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1429 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1428 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_INHSV3SR U1 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U4 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_XOR2HSV2 U6 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
endmodule


module cell_3_1427 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_46 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_46 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1457 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1456 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1455 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1454 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1453 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1452 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1451 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1450 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1449 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1448 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1447 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1446 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1445 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1444 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1443 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1442 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1441 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1440 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1439 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1438 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1437 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1436 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1435 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1434 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1433 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1432 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1431 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1430 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1429 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1428 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1427 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2 U1 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n2), .ZN(n3) );
  LVT_CLKNHSV0 U3 ( .I(t_m_1_in), .ZN(n2) );
endmodule


module cell_2_45 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_1426 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1425 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1424 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1423 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1422 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1421 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1420 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1419 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1418 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1417 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1416 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1415 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1414 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1413 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1412 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1411 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1410 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1409 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1408 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1407 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1406 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1405 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1404 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_NAND2HSV2 U1 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U3 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV0P5 U5 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_1403 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1402 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_1401 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1400 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1399 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_NAND2HSV2 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_NAND2HSV0P5 U4 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U5 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV2 U6 ( .I(n10), .ZN(n4) );
  LVT_INHSV0SR U7 ( .I(n9), .ZN(n5) );
  LVT_CLKNAND2HSV1 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_1398 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1397 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1396 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module row_other_45 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_45 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1426 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1425 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1424 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1423 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1422 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1421 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1420 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1419 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1418 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1417 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1416 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1415 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1414 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1413 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1412 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1411 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1410 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1409 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1408 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1407 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1406 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1405 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1404 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1403 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1402 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1401 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1400 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1399 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1398 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1397 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1396 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV6 U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_CLKNHSV16 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_44 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1395 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1394 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1393 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1392 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1391 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1390 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1389 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1388 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1387 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1386 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1385 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1384 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1383 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1382 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1381 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1380 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1379 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1378 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1377 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1376 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1375 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1374 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1373 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1372 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1371 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1370 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1369 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1368 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1367 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_XOR2HSV2 U1 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_CLKAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .Z(n3) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n3), .A2(t_i_1_in), .ZN(n4) );
endmodule


module cell_3_1366 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1365 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n6), .A2(n5), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2SR U4 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV2 U5 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U6 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV4 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_44 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_44 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1395 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1394 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1393 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1392 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1391 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1390 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1389 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1388 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1387 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1386 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1385 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1384 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1383 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1382 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1381 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1380 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1379 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1378 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1377 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1376 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1375 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1374 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1373 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1372 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1371 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1370 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1369 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1368 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1367 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1366 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1365 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV4SR U1 ( .I(t_m_1_in), .ZN(n2) );
  LVT_CLKNHSV4 U2 ( .I(n2), .ZN(n1) );
endmodule


module cell_2_43 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_1364 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1363 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1362 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1361 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1360 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1359 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1358 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1357 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1356 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1355 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1354 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1353 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1352 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1351 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1350 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1349 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1348 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1347 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1346 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1345 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1344 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1343 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1342 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1341 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1340 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1339 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1338 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1337 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1336 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_OAI21HSV2 U2 ( .A1(t_i_1_in), .A2(n5), .B(n2), .ZN(n4) );
  LVT_XNOR2HSV1 U3 ( .A1(n6), .A2(n4), .ZN(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(n5), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U5 ( .A1(b_in), .A2(a_in), .ZN(n5) );
endmodule


module cell_3_1335 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1334 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV4 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module row_other_43 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_43 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_1364 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1363 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1362 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1361 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1360 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1359 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1358 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1357 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1356 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1355 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1354 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1353 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1352 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1351 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1350 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1349 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1348 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1347 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1346 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1345 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1344 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1343 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1342 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1341 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1340 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1339 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1338 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1337 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1336 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1335 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1334 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV0SR U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_42 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_1333 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1332 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1331 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1330 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1329 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1328 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1327 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1326 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1325 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1324 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1323 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1322 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1321 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1320 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1319 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1318 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1317 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1316 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1315 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1314 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1313 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1312 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_1311 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_1310 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1309 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1308 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1307 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1306 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV3 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1305 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1304 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1303 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV3SR U1 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV0P5 U2 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U5 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_42 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_42 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1333 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1332 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1331 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1330 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1329 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1328 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1327 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1326 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1325 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1324 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1323 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1322 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1321 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1320 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1319 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1318 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1317 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1316 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1315 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1314 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1313 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1312 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1311 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1310 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1309 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1308 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1307 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1306 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1305 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1304 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1303 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV4 U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV8 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_41 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_1302 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1301 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1300 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1299 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1298 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1297 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1296 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1295 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1294 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1293 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1292 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1291 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1290 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1289 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1288 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1287 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1286 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1285 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1284 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1283 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1282 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1281 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1280 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1279 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1278 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1277 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U5 ( .I(n6), .ZN(n4) );
  LVT_XOR2HSV0 U6 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_3_1276 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1275 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV4 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_NAND2HSV1 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U5 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_3_1274 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1273 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_CLKNHSV2 U5 ( .I(n8), .ZN(n4) );
  LVT_XOR2HSV2 U6 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
endmodule


module cell_3_1272 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV4 U1 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_INHSV2 U6 ( .I(n10), .ZN(n4) );
  LVT_NAND2HSV0P5 U7 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_INHSV0SR U8 ( .I(n9), .ZN(n5) );
endmodule


module row_other_41 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_41 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1302 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1301 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1300 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1299 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1298 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1297 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1296 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1295 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1294 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1293 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1292 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1291 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1290 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1289 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1288 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1287 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1286 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1285 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1284 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1283 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1282 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1281 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1280 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1279 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1278 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1277 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1276 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1275 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1274 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1273 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1272 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV8 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV2SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_40 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_1271 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1270 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1269 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1268 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1267 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1266 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1265 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1264 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1263 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1262 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1261 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1260 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1259 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1258 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1257 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1256 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1255 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1254 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1253 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1252 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1251 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1250 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1249 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1248 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1247 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1246 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U4 ( .I(n6), .ZN(n4) );
  LVT_CLKXOR2HSV2 U5 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_1245 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1244 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1243 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1242 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_1241 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module row_other_40 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_40 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1271 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1270 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1269 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1268 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1267 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1266 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1265 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1264 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1263 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1262 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1261 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1260 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1259 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1258 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1257 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1256 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1255 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1254 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1253 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1252 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1251 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1250 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1249 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1248 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1247 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1246 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1245 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1244 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1243 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1242 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1241 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV8 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV2SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_39 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1240 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1239 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1238 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1237 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1236 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1235 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1234 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1233 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1232 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1231 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1230 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1229 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1228 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1227 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1226 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1225 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1224 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1223 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1222 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1221 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1220 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1219 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1218 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1217 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1216 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV1 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1215 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n2), .A2(n5), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_1214 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_1213 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1212 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1211 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1210 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_39 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_39 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1240 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1239 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1238 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1237 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1236 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1235 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1234 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1233 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1232 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1231 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1230 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1229 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1228 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1227 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1226 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1225 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1224 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1223 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1222 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1221 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1220 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1219 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1218 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1217 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1216 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1215 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1214 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1213 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1212 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1211 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1210 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV6 U1 ( .I(n3), .ZN(n1) );
  LVT_INHSV0P5 U2 ( .I(n3), .ZN(n2) );
  LVT_INHSV2SR U3 ( .I(t_m_1_in), .ZN(n3) );
endmodule


module cell_2_38 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1209 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1208 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1207 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1206 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1205 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1204 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1203 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1202 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1201 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1200 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1199 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1198 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1197 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1196 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1195 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1194 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1193 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1192 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1191 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1190 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1189 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1188 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1187 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1186 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1185 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1184 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1183 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1182 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1181 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1180 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1179 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XNOR2HSV4 U1 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNHSV4 U2 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV3 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV4 U6 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV4 U7 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNHSV4 U8 ( .I(n9), .ZN(n2) );
endmodule


module row_other_38 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_38 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_1209 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1208 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1207 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1206 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1205 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1204 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1203 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1202 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1201 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1200 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1199 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1198 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1197 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1196 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1195 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1194 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1193 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1192 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1191 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1190 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1189 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1188 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1187 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1186 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1185 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1184 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1183 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1182 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1181 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1180 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1179 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_37 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_1178 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1177 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1176 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1175 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1174 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1173 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1172 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1171 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1170 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1169 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1168 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1167 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1166 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1165 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1164 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1163 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1162 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1161 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1160 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1159 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1158 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1157 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1156 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1155 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1154 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1153 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1152 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1151 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1150 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1149 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1148 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U1 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV4 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNAND2HSV3 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNHSV2P5 U5 ( .I(n9), .ZN(n2) );
  LVT_XNOR2HSV4 U6 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
  LVT_CLKNAND2HSV3 U7 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U8 ( .I(n7), .ZN(n4) );
endmodule


module row_other_37 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_37 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_1178 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1177 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1176 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1175 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1174 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1173 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1172 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1171 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1170 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1169 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1168 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1167 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1166 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1165 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1164 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1163 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1162 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1161 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1160 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1159 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1158 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1157 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1156 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1155 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1154 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1153 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1152 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1151 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1150 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1149 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1148 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV4 U1 ( .I(n2), .ZN(n3) );
  LVT_INHSV3SR U2 ( .I(t_m_1_in), .ZN(n2) );
  LVT_CLKNHSV4 U3 ( .I(n2), .ZN(n1) );
endmodule


module cell_2_36 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1147 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1146 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1145 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1144 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n5), .A2(n6), .Z(t_i_out) );
endmodule


module cell_3_1143 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1142 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1141 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1140 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1139 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1138 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1137 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1136 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1135 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1134 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1133 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1132 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1131 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1130 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1129 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1128 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1127 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1126 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1125 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1124 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1123 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1122 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1121 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1120 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1119 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1118 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1117 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n6), .A2(n2), .ZN(n4) );
  LVT_CLKNAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U5 ( .A1(n8), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV2 U6 ( .I(t_i_1_in), .ZN(n2) );
  LVT_INHSV2 U7 ( .I(n8), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(n9), .A2(n7), .ZN(t_i_out) );
endmodule


module row_other_36 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_2_36 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1147 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1146 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1145 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1144 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1143 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1142 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1141 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1140 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1139 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1138 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1137 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1136 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1135 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1134 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1133 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1132 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1131 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1130 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1129 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1128 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1127 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1126 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1125 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1124 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1123 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1122 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1121 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1120 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1119 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1118 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1117 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2 U1 ( .I(t_m_1_in), .ZN(n3) );
  LVT_CLKNHSV4 U2 ( .I(n3), .ZN(n1) );
  LVT_CLKNHSV4 U3 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n4) );
endmodule


module cell_2_35 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1116 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1115 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1114 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1113 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1112 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_XOR2HSV0 U1 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_CLKNAND2HSV1 U3 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNAND2HSV3 U5 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_CLKNHSV0P5 U6 ( .I(n8), .ZN(n4) );
  LVT_CLKNHSV2P5 U7 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV8 U8 ( .A1(b_in), .A2(a_in), .ZN(n8) );
endmodule


module cell_3_1111 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1110 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1109 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1108 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1107 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1106 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1105 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1104 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1103 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1102 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1101 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1100 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1099 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1098 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1097 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1096 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1095 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1094 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1093 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1092 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV2 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U5 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0SR U6 ( .I(n8), .ZN(n4) );
  LVT_INHSV2 U7 ( .I(t_i_1_in), .ZN(n5) );
  LVT_CLKXOR2HSV2 U8 ( .A1(n10), .A2(n9), .Z(t_i_out) );
endmodule


module cell_3_1091 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1090 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1089 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1088 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n3, n4, n5;

  LVT_XOR2HSV2 U1 ( .A1(n5), .A2(n4), .Z(t_i_out) );
  LVT_XNOR2HSV1 U2 ( .A1(n3), .A2(t_i_1_in), .ZN(n4) );
  LVT_CLKAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .Z(n3) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_1087 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV2 U4 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
endmodule


module cell_3_1086 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_INHSV2SR U1 ( .I(n9), .ZN(n2) );
  LVT_CLKNAND2HSV1 U2 ( .A1(n9), .A2(n7), .ZN(n6) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n2), .A2(n4), .ZN(n5) );
  LVT_CLKNAND2HSV3 U5 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNHSV2 U6 ( .I(n7), .ZN(n4) );
  LVT_CLKNAND2HSV2 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV4 U8 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
endmodule


module row_other_35 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_2_35 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_1116 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1115 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1114 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1113 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1112 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1111 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1110 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1109 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1108 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1107 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1106 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1105 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1104 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1103 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1102 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1101 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1100 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1099 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1098 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1097 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1096 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1095 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1094 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1093 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1092 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1091 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1090 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n4), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1089 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1088 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1087 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1086 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV2 U1 ( .I(t_m_1_in), .ZN(n3) );
  LVT_CLKNHSV8 U2 ( .I(n3), .ZN(n4) );
  LVT_INHSV0SR U3 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_34 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_1085 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1084 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1083 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_XOR2HSV0 U1 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U2 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U5 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0SR U6 ( .I(n8), .ZN(n4) );
  LVT_INHSV2 U7 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV2 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_1082 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1081 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1080 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1079 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1078 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1077 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1076 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1075 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1074 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1073 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
endmodule


module cell_3_1072 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1071 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0SR U5 ( .I(n8), .ZN(n4) );
  LVT_INHSV2 U6 ( .I(t_i_1_in), .ZN(n5) );
  LVT_XOR2HSV4 U7 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_1070 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1069 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1068 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1067 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1066 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1065 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1064 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1063 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1062 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1061 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1060 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1059 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1058 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1057 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1056 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1055 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n2), .A2(n4), .ZN(n5) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNHSV2P5 U4 ( .I(n9), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV3 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV1 U7 ( .A1(n9), .A2(n7), .ZN(n6) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_34 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_34 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_1085 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1084 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1083 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1082 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1081 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1080 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1079 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1078 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1077 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1076 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1075 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1074 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1073 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1072 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1071 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1070 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1069 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1068 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1067 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1066 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1065 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1064 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1063 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1062 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1061 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1060 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1059 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1058 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n3), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1057 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1056 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1055 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV3SR U1 ( .I(n2), .ZN(n1) );
  LVT_INHSV2SR U2 ( .I(t_m_1_in), .ZN(n2) );
  LVT_INHSV4 U3 ( .I(n2), .ZN(n3) );
endmodule


module cell_2_33 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1054 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1053 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1052 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1051 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1050 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1049 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1048 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1047 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1046 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1045 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1044 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1043 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1042 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1041 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1040 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1039 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1038 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1037 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1036 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1035 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1034 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1033 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1032 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1031 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1030 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1029 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1028 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1027 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1026 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1025 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_CLKNAND2HSV2 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0P5 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNAND2HSV3 U3 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_CLKNHSV0 U5 ( .I(n8), .ZN(n4) );
  LVT_CLKNHSV2 U6 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV0 U7 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV2 U8 ( .A1(n10), .A2(n9), .Z(t_i_out) );
endmodule


module cell_3_1024 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_INAND2HSV4 U1 ( .A1(n9), .B1(n8), .ZN(n6) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XOR2HSV2 U5 ( .A1(n7), .A2(t_i_1_in), .Z(n8) );
  LVT_INHSV2SR U6 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0P5 U7 ( .A1(n9), .A2(n4), .ZN(n5) );
endmodule


module row_other_33 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_33 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_1054 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1053 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1052 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1051 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1050 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1049 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1048 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1047 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1046 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1045 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1044 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1043 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1042 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1041 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1040 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1039 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1038 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1037 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1036 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1035 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1034 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1033 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1032 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1031 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_1030 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_1029 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_1028 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_1027 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_1026 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        n1), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1025 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_1024 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV8RT U1 ( .I(t_m_1_in), .Z(n1) );
  LVT_INHSV2 U2 ( .I(n2), .ZN(n3) );
  LVT_INHSV0SR U3 ( .I(t_m_1_in), .ZN(n2) );
endmodule


module cell_2_32 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_1023 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1022 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1021 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1020 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1019 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1018 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1017 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0P5 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_CLKNHSV0P5 U5 ( .I(n10), .ZN(n4) );
  LVT_CLKNHSV0P5 U6 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV0 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_XOR2HSV2 U8 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
endmodule


module cell_3_1016 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1015 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1014 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1013 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1012 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1011 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_1010 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0P5 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_CLKNHSV0P5 U5 ( .I(n10), .ZN(n4) );
  LVT_INHSV2SR U6 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV0 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_XOR2HSV2 U8 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
endmodule


module cell_3_1009 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1008 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1007 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1006 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV2 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_CLKNAND2HSV1 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNAND2HSV2 U5 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_CLKNHSV0 U6 ( .I(n8), .ZN(n4) );
  LVT_INHSV2 U7 ( .I(t_i_1_in), .ZN(n5) );
  LVT_XOR2HSV2 U8 ( .A1(n10), .A2(n9), .Z(t_i_out) );
endmodule


module cell_3_1005 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1004 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1003 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1002 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1001 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_1000 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_999 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_998 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_997 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_996 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_995 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_994 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_993 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_32 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_32 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_1023 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_1022 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_1021 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_1020 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_1019 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_1018 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_1017 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_1016 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_1015 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_1014 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_1013 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_1012 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_1011 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_1010 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_1009 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_1008 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_1007 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_1006 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_1005 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_1004 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_1003 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_1002 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_1001 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_1000 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_999 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_998 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_997 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_996 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_995 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_994 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_993 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_31 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n3), .A2(n4), .Z(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_992 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV1 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_991 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_990 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV1 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_989 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_OAI21HSV0 U1 ( .A1(n6), .A2(n4), .B(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(n6), .A2(n4), .ZN(n2) );
  LVT_XNOR2HSV1 U4 ( .A1(n5), .A2(t_i_1_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_988 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_OAI21HSV0 U1 ( .A1(n6), .A2(n4), .B(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U2 ( .A1(n6), .A2(n4), .ZN(n2) );
  LVT_XNOR2HSV1 U4 ( .A1(n5), .A2(t_i_1_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_987 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV1 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_986 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_985 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_984 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_983 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_982 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_981 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_980 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV2 U5 ( .I(n8), .ZN(n4) );
  LVT_INHSV2 U6 ( .I(t_i_1_in), .ZN(n5) );
  LVT_XOR2HSV0 U7 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_979 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_978 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_977 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_976 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_975 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_974 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_973 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0SR U5 ( .I(n8), .ZN(n4) );
  LVT_INHSV2 U6 ( .I(t_i_1_in), .ZN(n5) );
  LVT_XOR2HSV0 U7 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_972 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_971 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_970 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_969 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_968 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0SR U5 ( .I(n8), .ZN(n4) );
  LVT_INHSV2SR U6 ( .I(t_i_1_in), .ZN(n5) );
  LVT_XOR2HSV0 U7 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_967 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_966 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_965 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_964 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_XNOR2HSV1 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_963 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_962 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module row_other_31 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_31 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_992 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_991 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_990 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_989 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_988 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_987 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_986 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_985 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_984 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_983 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_982 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_981 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_980 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_979 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_978 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_977 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_976 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_975 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_974 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_973 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_972 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_971 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_970 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_969 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_968 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_967 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_966 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_965 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_964 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_963 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_962 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_1 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [31:0] a_in;
  input [31:0] g_in;
  input [31:0] b_in;
  input [31:0] t_m_1_in;
  input [30:0] t_i_1_in;
  input [30:0] t_i_2_in;
  output [31:0] a_out;
  output [31:0] g_out;
  output [30:0] t_i_1_out;
  output [30:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;
  wire   n1, n2, n4, n5, n7, n8, n10, n12, n14, n15;
  wire   [30:0] t0;
  wire   [30:0] t1;
  wire   [30:0] t2;
  wire   [30:0] t3;
  wire   [30:0] t4;
  wire   [30:0] t5;
  wire   [30:0] t6;
  wire   [30:0] t7;
  wire   [30:0] t8;
  wire   [30:0] t9;
  wire   [30:0] t10;
  wire   [30:0] t11;
  wire   [30:0] t12;
  wire   [30:0] t13;
  wire   [30:0] t14;
  wire   [30:0] t15;
  wire   [30:0] t16;
  wire   [30:0] t17;
  wire   [30:0] t18;
  wire   [30:0] t19;
  wire   [30:0] t20;
  wire   [30:0] t21;
  wire   [30:0] t22;
  wire   [30:0] t23;
  wire   [30:0] t24;
  wire   [30:0] t25;
  wire   [30:0] t26;
  wire   [30:0] t27;
  wire   [30:0] t28;
  wire   [30:0] t29;
  wire   [30:0] t30;
  assign a_out[30] = a_in[30];
  assign a_out[29] = a_in[29];
  assign a_out[28] = a_in[28];
  assign a_out[27] = a_in[27];
  assign a_out[26] = a_in[26];
  assign a_out[25] = a_in[25];
  assign a_out[24] = a_in[24];
  assign a_out[23] = a_in[23];
  assign a_out[22] = a_in[22];
  assign a_out[20] = a_in[20];
  assign a_out[19] = a_in[19];
  assign a_out[18] = a_in[18];
  assign a_out[17] = a_in[17];
  assign a_out[16] = a_in[16];
  assign a_out[15] = a_in[15];
  assign a_out[14] = a_in[14];
  assign a_out[13] = a_in[13];
  assign a_out[12] = a_in[12];
  assign a_out[11] = a_in[11];
  assign a_out[10] = a_in[10];
  assign a_out[9] = a_in[9];
  assign a_out[8] = a_in[8];
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[29] = g_in[29];
  assign g_out[28] = g_in[28];
  assign g_out[27] = g_in[27];
  assign g_out[26] = g_in[26];
  assign g_out[25] = g_in[25];
  assign g_out[24] = g_in[24];
  assign g_out[23] = g_in[23];
  assign g_out[22] = g_in[22];
  assign g_out[20] = g_in[20];
  assign g_out[19] = g_in[19];
  assign g_out[18] = g_in[18];
  assign g_out[17] = g_in[17];
  assign g_out[16] = g_in[16];
  assign g_out[15] = g_in[15];
  assign g_out[14] = g_in[14];
  assign g_out[13] = g_in[13];
  assign g_out[12] = g_in[12];
  assign g_out[11] = g_in[11];
  assign g_out[10] = g_in[10];
  assign g_out[9] = g_in[9];
  assign g_out[8] = g_in[8];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_1 u0 ( .a_in({a_in[31:22], n8, a_in[20:0]}), .g_in({g_in[31], n2, 
        g_in[29:22], n5, g_in[20:0]}), .b_in(b_in[31]), .t_m_1_in(t_m_1_in[31]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), .t_i_2_in(t_i_2_in), .t_i_1_out(t0), 
        .t_i_2_out(t_i_2_out[30]) );
  row_other_61 u1 ( .a_in({a_in[31:22], a_out[21], a_in[20:0]}), .g_in({
        g_in[31], g_out[30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[30]), .t_m_1_in(t_m_1_in[30]), .t_i_1_in(t0), .t_i_1_out(t1), 
        .t_i_2_out(t_i_2_out[29]) );
  row_other_60 u2 ( .a_in({a_in[31:22], a_out[21], a_in[20:0]}), .g_in({
        g_in[31], g_out[30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[29]), .t_m_1_in(t_m_1_in[29]), .t_i_1_in(t1), .t_i_1_out(t2), 
        .t_i_2_out(t_i_2_out[28]) );
  row_other_59 u3 ( .a_in({a_in[31:22], a_out[21], a_in[20:0]}), .g_in({
        g_in[31], g_out[30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[28]), .t_m_1_in(t_m_1_in[28]), .t_i_1_in(t2), .t_i_1_out(t3), 
        .t_i_2_out(t_i_2_out[27]) );
  row_other_58 u4 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_in[31], g_out[30], g_in[29:22], g_out[21], g_in[20:0]}), 
        .b_in(b_in[27]), .t_m_1_in(t_m_1_in[27]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(t_i_2_out[26]) );
  row_other_57 u5 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_in[31], g_out[30], g_in[29:22], g_out[21], g_in[20:0]}), 
        .b_in(b_in[26]), .t_m_1_in(t_m_1_in[26]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(t_i_2_out[25]) );
  row_other_56 u6 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_in[31], g_out[30], g_in[29:22], g_out[21], g_in[20:0]}), 
        .b_in(b_in[25]), .t_m_1_in(t_m_1_in[25]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(t_i_2_out[24]) );
  row_other_55 u7 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_in[31], g_out[30], g_in[29:22], g_out[21], g_in[20:0]}), 
        .b_in(b_in[24]), .t_m_1_in(t_m_1_in[24]), .t_i_1_in(t6), .t_i_1_out(t7), .t_i_2_out(t_i_2_out[23]) );
  row_other_54 u8 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[23]), .t_m_1_in(t_m_1_in[23]), .t_i_1_in(t7), .t_i_1_out(t8), 
        .t_i_2_out(t_i_2_out[22]) );
  row_other_53 u9 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[22]), .t_m_1_in(t_m_1_in[22]), .t_i_1_in(t8), .t_i_1_out(t9), 
        .t_i_2_out(t_i_2_out[21]) );
  row_other_52 u10 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[21]), .t_m_1_in(t_m_1_in[21]), .t_i_1_in(t9), .t_i_1_out(t10), 
        .t_i_2_out(t_i_2_out[20]) );
  row_other_51 u11 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[20]), .t_m_1_in(t_m_1_in[20]), .t_i_1_in(t10), .t_i_1_out(t11), 
        .t_i_2_out(t_i_2_out[19]) );
  row_other_50 u12 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[19]), .t_m_1_in(t_m_1_in[19]), .t_i_1_in(t11), .t_i_1_out(t12), 
        .t_i_2_out(t_i_2_out[18]) );
  row_other_49 u13 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[18]), .t_m_1_in(t_m_1_in[18]), .t_i_1_in(t12), .t_i_1_out(t13), 
        .t_i_2_out(t_i_2_out[17]) );
  row_other_48 u14 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[17]), .t_m_1_in(t_m_1_in[17]), .t_i_1_in(t13), .t_i_1_out(t14), 
        .t_i_2_out(t_i_2_out[16]) );
  row_other_47 u15 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[16]), .t_m_1_in(t_m_1_in[16]), .t_i_1_in(t14), .t_i_1_out(t15), 
        .t_i_2_out(t_i_2_out[15]) );
  row_other_46 u16 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[15]), .t_m_1_in(t_m_1_in[15]), .t_i_1_in(t15), .t_i_1_out(t16), 
        .t_i_2_out(t_i_2_out[14]) );
  row_other_45 u17 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[14]), .t_m_1_in(t_m_1_in[14]), .t_i_1_in(t16), .t_i_1_out(t17), 
        .t_i_2_out(t_i_2_out[13]) );
  row_other_44 u18 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[13]), .t_m_1_in(t_m_1_in[13]), .t_i_1_in(t17), .t_i_1_out(t18), 
        .t_i_2_out(t_i_2_out[12]) );
  row_other_43 u19 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[12]), .t_m_1_in(t_m_1_in[12]), .t_i_1_in(t18), .t_i_1_out(t19), 
        .t_i_2_out(t_i_2_out[11]) );
  row_other_42 u20 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[11]), .t_m_1_in(t_m_1_in[11]), .t_i_1_in(t19), .t_i_1_out(t20), 
        .t_i_2_out(t_i_2_out[10]) );
  row_other_41 u21 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[10]), .t_m_1_in(t_m_1_in[10]), .t_i_1_in(t20), .t_i_1_out(t21), 
        .t_i_2_out(t_i_2_out[9]) );
  row_other_40 u22 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[9]), .t_m_1_in(t_m_1_in[9]), .t_i_1_in(t21), .t_i_1_out(t22), 
        .t_i_2_out(t_i_2_out[8]) );
  row_other_39 u23 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[8]), .t_m_1_in(t_m_1_in[8]), .t_i_1_in(t22), .t_i_1_out(t23), 
        .t_i_2_out(t_i_2_out[7]) );
  row_other_38 u24 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[7]), .t_m_1_in(n15), .t_i_1_in(t23), .t_i_1_out(t24), .t_i_2_out(
        t_i_2_out[6]) );
  row_other_37 u25 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[6]), .t_m_1_in(t_m_1_in[6]), .t_i_1_in(t24), .t_i_1_out(t25), 
        .t_i_2_out(t_i_2_out[5]) );
  row_other_36 u26 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[5]), .t_m_1_in(t_m_1_in[5]), .t_i_1_in(t25), .t_i_1_out(t26), 
        .t_i_2_out(t_i_2_out[4]) );
  row_other_35 u27 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[4]), .t_m_1_in(t_m_1_in[4]), .t_i_1_in(t26), .t_i_1_out(t27), 
        .t_i_2_out(t_i_2_out[3]) );
  row_other_34 u28 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[3]), .t_m_1_in(t_m_1_in[3]), .t_i_1_in(t27), .t_i_1_out(t28), 
        .t_i_2_out(t_i_2_out[2]) );
  row_other_33 u29 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[2]), .t_m_1_in(t_m_1_in[2]), .t_i_1_in(t28), .t_i_1_out(t29), 
        .t_i_2_out(t_i_2_out[1]) );
  row_other_32 u30 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[1]), .t_m_1_in(t_m_1_in[1]), .t_i_1_in(t29), .t_i_1_out(t30), 
        .t_i_2_out(t_i_2_out[0]) );
  row_other_31 u31 ( .a_in({a_out[31], a_in[30:22], a_out[21], a_in[20:0]}), 
        .g_in({g_out[31:30], g_in[29:22], g_out[21], g_in[20:0]}), .b_in(
        b_in[0]), .t_m_1_in(t_m_1_in[0]), .t_i_1_in(t30), .t_i_1_out(t_i_1_out), .t_i_2_out(t_i_1_out_0) );
  LVT_INHSV8SR U1 ( .I(t_m_1_in[7]), .ZN(n14) );
  LVT_CLKNHSV16 U2 ( .I(n14), .ZN(n15) );
  LVT_INHSV4 U3 ( .I(g_in[30]), .ZN(n1) );
  LVT_INHSV2P5 U4 ( .I(n1), .ZN(n2) );
  LVT_INHSV2SR U5 ( .I(n1), .ZN(g_out[30]) );
  LVT_INHSV2 U6 ( .I(n4), .ZN(n5) );
  LVT_INHSV2 U7 ( .I(a_in[21]), .ZN(n7) );
  LVT_INHSV2 U8 ( .I(g_in[21]), .ZN(n4) );
  LVT_INHSV2SR U9 ( .I(n4), .ZN(g_out[21]) );
  LVT_CLKNHSV2 U10 ( .I(n7), .ZN(n8) );
  LVT_INHSV2SR U11 ( .I(n7), .ZN(a_out[21]) );
  LVT_INHSV0SR U12 ( .I(a_in[31]), .ZN(n10) );
  LVT_INHSV2 U13 ( .I(n10), .ZN(a_out[31]) );
  LVT_INHSV0SR U14 ( .I(g_in[31]), .ZN(n12) );
  LVT_CLKNHSV4 U15 ( .I(n12), .ZN(g_out[31]) );
endmodule


module regist_32bit_7 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_32bit_6 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_31bit_4 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n2), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n2), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module PE_1 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro );
  input [31:0] a_in;
  input [31:0] g_in;
  input [31:0] b_in;
  input [30:0] t_i_1_in;
  input [30:0] t_i_2_in;
  output [31:0] a_out;
  output [31:0] g_out;
  output [31:0] b_out;
  output [30:0] t_i_1_out;
  output [30:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   n104, n105, n106, l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0,
         to_1, ti_1, n14, n15, n16, n17, n18, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103;
  wire   [31:0] l_a;
  wire   [31:0] l_g;
  wire   [30:0] l_t_i_1_in;
  wire   [30:0] l_t_i_2_in;
  wire   [31:0] mux_b;
  wire   [31:0] mux_bq;
  wire   [30:0] to_7;
  wire   [30:0] ti_7;
  wire   [31:0] ao;
  wire   [31:0] go;
  wire   [30:0] to;

  LVT_AO22HSV0 U35 ( .A1(mux_bq[9]), .A2(n83), .B1(b_out[9]), .B2(n90), .Z(
        mux_b[9]) );
  LVT_AO22HSV0 U36 ( .A1(mux_bq[8]), .A2(n83), .B1(b_out[8]), .B2(n90), .Z(
        mux_b[8]) );
  LVT_AO22HSV0 U37 ( .A1(mux_bq[7]), .A2(n83), .B1(b_out[7]), .B2(n90), .Z(
        mux_b[7]) );
  LVT_AO22HSV0 U38 ( .A1(mux_bq[6]), .A2(n83), .B1(b_out[6]), .B2(n90), .Z(
        mux_b[6]) );
  LVT_AO22HSV0 U39 ( .A1(mux_bq[5]), .A2(n83), .B1(b_out[5]), .B2(n90), .Z(
        mux_b[5]) );
  LVT_AO22HSV0 U40 ( .A1(mux_bq[4]), .A2(n83), .B1(b_out[4]), .B2(n90), .Z(
        mux_b[4]) );
  LVT_AO22HSV0 U41 ( .A1(mux_bq[3]), .A2(n83), .B1(b_out[3]), .B2(n90), .Z(
        mux_b[3]) );
  LVT_AO22HSV0 U44 ( .A1(mux_bq[2]), .A2(n83), .B1(b_out[2]), .B2(n90), .Z(
        mux_b[2]) );
  LVT_AO22HSV0 U47 ( .A1(mux_bq[27]), .A2(n83), .B1(b_out[27]), .B2(n90), .Z(
        mux_b[27]) );
  LVT_AO22HSV0 U48 ( .A1(mux_bq[26]), .A2(n83), .B1(b_out[26]), .B2(n90), .Z(
        mux_b[26]) );
  LVT_AO22HSV0 U49 ( .A1(mux_bq[25]), .A2(n83), .B1(b_out[25]), .B2(n90), .Z(
        mux_b[25]) );
  LVT_AO22HSV0 U50 ( .A1(mux_bq[24]), .A2(n83), .B1(b_out[24]), .B2(n90), .Z(
        mux_b[24]) );
  LVT_AO22HSV0 U51 ( .A1(mux_bq[23]), .A2(n83), .B1(b_out[23]), .B2(n90), .Z(
        mux_b[23]) );
  LVT_AO22HSV0 U52 ( .A1(mux_bq[22]), .A2(n83), .B1(b_out[22]), .B2(n90), .Z(
        mux_b[22]) );
  LVT_AO22HSV0 U53 ( .A1(mux_bq[21]), .A2(n83), .B1(b_out[21]), .B2(n90), .Z(
        mux_b[21]) );
  LVT_AO22HSV0 U54 ( .A1(mux_bq[20]), .A2(n83), .B1(b_out[20]), .B2(n90), .Z(
        mux_b[20]) );
  LVT_AO22HSV0 U55 ( .A1(mux_bq[1]), .A2(n83), .B1(b_out[1]), .B2(n90), .Z(
        mux_b[1]) );
  LVT_AO22HSV0 U56 ( .A1(mux_bq[19]), .A2(n83), .B1(b_out[19]), .B2(n90), .Z(
        mux_b[19]) );
  LVT_AO22HSV0 U57 ( .A1(mux_bq[18]), .A2(n83), .B1(b_out[18]), .B2(n90), .Z(
        mux_b[18]) );
  LVT_AO22HSV0 U58 ( .A1(mux_bq[17]), .A2(n83), .B1(b_out[17]), .B2(n90), .Z(
        mux_b[17]) );
  LVT_AO22HSV0 U59 ( .A1(mux_bq[16]), .A2(n83), .B1(b_out[16]), .B2(n90), .Z(
        mux_b[16]) );
  LVT_AO22HSV0 U60 ( .A1(mux_bq[15]), .A2(n83), .B1(b_out[15]), .B2(n90), .Z(
        mux_b[15]) );
  LVT_AO22HSV0 U61 ( .A1(mux_bq[14]), .A2(n83), .B1(b_out[14]), .B2(n90), .Z(
        mux_b[14]) );
  LVT_AO22HSV0 U62 ( .A1(mux_bq[13]), .A2(n83), .B1(b_out[13]), .B2(n90), .Z(
        mux_b[13]) );
  LVT_AO22HSV0 U63 ( .A1(mux_bq[12]), .A2(n83), .B1(b_out[12]), .B2(n90), .Z(
        mux_b[12]) );
  LVT_AO22HSV0 U64 ( .A1(mux_bq[11]), .A2(n83), .B1(b_out[11]), .B2(n90), .Z(
        mux_b[11]) );
  LVT_AO22HSV0 U65 ( .A1(mux_bq[10]), .A2(n83), .B1(b_out[10]), .B2(n90), .Z(
        mux_b[10]) );
  LVT_AO22HSV0 U66 ( .A1(mux_bq[0]), .A2(n83), .B1(b_out[0]), .B2(n90), .Z(
        mux_b[0]) );
  LVT_NOR2HSV0 U67 ( .A1(n102), .A2(n90), .ZN(c_t_i_1_in_0) );
  LVT_AOI21HSV0 U69 ( .A1(n100), .A2(n99), .B(n90), .ZN(\c_t_i_1_in[0] ) );
  LVT_AND4HSV0 U71 ( .A1(n98), .A2(n97), .A3(n96), .A4(n95), .Z(n99) );
  LVT_NOR4HSV0 U72 ( .A1(l_t_i_1_in[9]), .A2(l_t_i_1_in[8]), .A3(l_t_i_1_in[7]), .A4(l_t_i_1_in[6]), .ZN(n95) );
  LVT_NOR4HSV0 U73 ( .A1(l_t_i_1_in[5]), .A2(l_t_i_1_in[4]), .A3(l_t_i_1_in[3]), .A4(l_t_i_1_in[30]), .ZN(n96) );
  LVT_NOR4HSV0 U74 ( .A1(l_t_i_1_in[2]), .A2(l_t_i_1_in[29]), .A3(
        l_t_i_1_in[28]), .A4(l_t_i_1_in[27]), .ZN(n97) );
  LVT_NOR4HSV0 U75 ( .A1(l_t_i_1_in[26]), .A2(l_t_i_1_in[25]), .A3(
        l_t_i_1_in[24]), .A4(l_t_i_1_in[23]), .ZN(n98) );
  LVT_AND4HSV0 U76 ( .A1(n94), .A2(n93), .A3(n92), .A4(n91), .Z(n100) );
  LVT_NOR4HSV0 U77 ( .A1(l_t_i_1_in[22]), .A2(l_t_i_1_in[21]), .A3(
        l_t_i_1_in[20]), .A4(l_t_i_1_in[1]), .ZN(n91) );
  LVT_NOR4HSV0 U78 ( .A1(l_t_i_1_in[19]), .A2(l_t_i_1_in[18]), .A3(
        l_t_i_1_in[17]), .A4(l_t_i_1_in[16]), .ZN(n92) );
  LVT_NOR4HSV0 U79 ( .A1(l_t_i_1_in[15]), .A2(l_t_i_1_in[14]), .A3(
        l_t_i_1_in[13]), .A4(l_t_i_1_in[12]), .ZN(n93) );
  LVT_NOR3HSV0 U80 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[11]), .A3(
        l_t_i_1_in[10]), .ZN(n94) );
  regist_32bit_11 u0 ( .clk(clk), .rstn(rstn), .in(a_in), .out(l_a) );
  regist_32bit_10 u1 ( .clk(clk), .rstn(rstn), .in(b_in), .out(b_out) );
  regist_32bit_9 u2 ( .clk(clk), .rstn(rstn), .in(g_in), .out(l_g) );
  regist_1bit_7 u3 ( .clk(clk), .rstn(rstn), .in(ctr), .out(l_ctr) );
  regist_1bit_6 u4 ( .clk(clk), .rstn(rstn), .in(n83), .out(n106) );
  regist_31bit_7 u5 ( .clk(clk), .rstn(rstn), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_31bit_6 u6 ( .clk(clk), .rstn(rstn), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_5 u7 ( .clk(clk), .rstn(rstn), .in(t_i_1_in_0), .out(
        l_t_i_1_in_0) );
  regist_32bit_8 u9 ( .clk(clk), .rstn(rstn), .in(mux_b), .out(mux_bq) );
  regist_1bit_4 u10 ( .clk(clk), .rstn(rstn), .in(to_1), .out(ti_1) );
  regist_31bit_5 u11 ( .clk(clk), .rstn(rstn), .in({to_7[30], n73, n63, 
        to_7[27:25], n31, n74, to_7[22:20], n72, to_7[18:17], n49, to_7[15:14], 
        n80, to_7[12], n81, n82, n75, to_7[8:5], n46, n76, n77, n78, n79}), 
        .out(ti_7) );
  PE_core_1 pe ( .a_in(l_a), .g_in(l_g), .b_in({n29, mux_bq[30:0]}), 
        .t_m_1_in({to_1, to_7[30], n73, n63, to_7[27:25], n31, n74, 
        to_7[22:17], n49, to_7[15:14], n80, to_7[12], n81, n82, n75, to_7[8:4], 
        n76, n77, n78, n79}), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \c_t_i_1_in[0] }), .t_i_1_in_0(c_t_i_1_in_0), .t_i_2_in(l_t_i_2_in), 
        .a_out(ao), .g_out(go), .t_i_1_out(to), .t_i_2_out({t_i_2_out[30:18], 
        n104, t_i_2_out[16:8], n105, t_i_2_out[6:0]}), .t_i_1_out_0(
        t_i_1_out_0) );
  regist_32bit_7 u12 ( .clk(clk), .rstn(rstn), .in(ao), .out(a_out) );
  regist_32bit_6 u13 ( .clk(clk), .rstn(rstn), .in(go), .out(g_out) );
  regist_31bit_4 u14 ( .clk(clk), .rstn(rstn), .in(to), .out(t_i_1_out) );
  LVT_NAND2HSV8 U2 ( .A1(n85), .A2(n84), .ZN(to_7[14]) );
  LVT_INHSV10SR U3 ( .I(n62), .ZN(n79) );
  LVT_AO22HSV2 U4 ( .A1(ti_7[20]), .A2(ctro), .B1(t_i_2_out[20]), .B2(n16), 
        .Z(to_7[20]) );
  LVT_NAND2HSV4 U5 ( .A1(n26), .A2(n27), .ZN(to_7[17]) );
  LVT_INHSV6 U6 ( .I(n59), .ZN(n76) );
  LVT_CLKNHSV6 U7 ( .I(n42), .ZN(n73) );
  LVT_NAND2HSV4 U8 ( .A1(n104), .A2(n16), .ZN(n27) );
  LVT_CLKNHSV2P5 U9 ( .I(n38), .ZN(n74) );
  LVT_AND2HSV4 U10 ( .A1(t_i_2_out[27]), .A2(n16), .Z(n57) );
  LVT_INHSV3SR U11 ( .I(n39), .ZN(n49) );
  LVT_INHSV6 U12 ( .I(n58), .ZN(n63) );
  LVT_CLKNAND2HSV3 U13 ( .A1(t_i_2_out[5]), .A2(n16), .ZN(n37) );
  LVT_INHSV10 U14 ( .I(n30), .ZN(n31) );
  LVT_INHSV4 U15 ( .I(n17), .ZN(n30) );
  LVT_OR2HSV4RQ U16 ( .A1(n51), .A2(n50), .Z(n72) );
  LVT_INHSV4SR U17 ( .I(n32), .ZN(n82) );
  LVT_NAND2HSV4 U18 ( .A1(n24), .A2(n25), .ZN(to_7[22]) );
  LVT_INHSV10 U19 ( .I(n35), .ZN(n78) );
  LVT_OR2HSV12RD U20 ( .A1(n67), .A2(n66), .Z(to_7[18]) );
  LVT_AND2HSV4 U21 ( .A1(t_i_2_out[18]), .A2(n16), .Z(n67) );
  LVT_CLKNAND2HSV3 U22 ( .A1(ti_1), .A2(l_ctr), .ZN(n88) );
  LVT_NAND2HSV4 U23 ( .A1(n37), .A2(n36), .ZN(to_7[5]) );
  LVT_INHSV4SR U24 ( .I(n103), .ZN(n14) );
  LVT_CLKNHSV2P5 U25 ( .I(n14), .ZN(n15) );
  LVT_INHSV4SR U26 ( .I(n14), .ZN(n16) );
  LVT_OR2HSV12RD U27 ( .A1(n51), .A2(n50), .Z(to_7[19]) );
  LVT_AOI22HSV2 U28 ( .A1(ti_7[23]), .A2(ctro), .B1(t_i_2_out[23]), .B2(n16), 
        .ZN(n38) );
  LVT_CLKAND2HSV4 U29 ( .A1(t_i_2_out[19]), .A2(n16), .Z(n51) );
  LVT_CLKNHSV4 U30 ( .I(n18), .ZN(n103) );
  LVT_NAND2HSV2 U31 ( .A1(t_i_2_out[8]), .A2(n16), .ZN(n53) );
  LVT_NAND2HSV2 U32 ( .A1(n22), .A2(n23), .ZN(n17) );
  LVT_INHSV8 U33 ( .I(n60), .ZN(n77) );
  LVT_CLKNHSV10 U34 ( .I(l_ctr), .ZN(n101) );
  LVT_OR2HSV12RD U42 ( .A1(n57), .A2(n56), .Z(to_7[27]) );
  LVT_BUFHSV2 U43 ( .I(n106), .Z(n18) );
  LVT_BUFHSV4 U45 ( .I(n106), .Z(ctro) );
  LVT_AND2HSV4 U46 ( .A1(t_i_2_out[10]), .A2(n16), .Z(n21) );
  LVT_INHSV4SR U68 ( .I(n41), .ZN(n75) );
  LVT_INHSV4SR U70 ( .I(n40), .ZN(n80) );
  LVT_CLKNAND2HSV4 U81 ( .A1(n69), .A2(n68), .ZN(to_7[26]) );
  LVT_NAND2HSV4 U82 ( .A1(t_i_2_out[22]), .A2(n16), .ZN(n25) );
  LVT_CLKNAND2HSV4 U83 ( .A1(n65), .A2(n64), .ZN(to_7[4]) );
  LVT_NAND2HSV4 U84 ( .A1(t_i_2_out[4]), .A2(n16), .ZN(n65) );
  LVT_NAND2HSV4 U85 ( .A1(n52), .A2(n53), .ZN(to_7[8]) );
  LVT_NAND2HSV2 U86 ( .A1(ti_7[24]), .A2(ctro), .ZN(n22) );
  LVT_CLKNHSV16 U87 ( .I(n28), .ZN(n29) );
  LVT_CLKNHSV8 U88 ( .I(mux_bq[31]), .ZN(n28) );
  LVT_NAND2HSV0P5 U89 ( .A1(t_i_2_out[24]), .A2(n16), .ZN(n23) );
  LVT_NAND2HSV4 U90 ( .A1(t_i_2_out[14]), .A2(n16), .ZN(n85) );
  LVT_CLKNAND2HSV8 U91 ( .A1(n88), .A2(n89), .ZN(to_1) );
  LVT_NAND2HSV4 U92 ( .A1(t_i_2_out[26]), .A2(n16), .ZN(n69) );
  LVT_NAND2HSV8 U93 ( .A1(n71), .A2(n70), .ZN(to_7[6]) );
  LVT_NAND2HSV4 U94 ( .A1(t_i_2_out[6]), .A2(n16), .ZN(n71) );
  LVT_AND2HSV2RD U95 ( .A1(ti_7[10]), .A2(ctro), .Z(n20) );
  LVT_NOR2HSV4 U96 ( .A1(n20), .A2(n21), .ZN(n32) );
  LVT_CLKNAND2HSV1 U97 ( .A1(ti_7[22]), .A2(ctro), .ZN(n24) );
  LVT_NAND2HSV2 U98 ( .A1(ti_7[17]), .A2(ctro), .ZN(n26) );
  LVT_INHSV2 U99 ( .I(ti_7[7]), .ZN(n34) );
  LVT_OR2HSV12RD U100 ( .A1(n48), .A2(n47), .Z(to_7[15]) );
  LVT_OR2HSV12RD U101 ( .A1(n55), .A2(n54), .Z(to_7[12]) );
  LVT_INHSV2 U102 ( .I(n33), .ZN(n90) );
  LVT_INHSV0SR U103 ( .I(n101), .ZN(n33) );
  LVT_INHSV4SR U104 ( .I(n61), .ZN(n81) );
  LVT_MOAI22HSV4 U105 ( .A1(n34), .A2(n16), .B1(n105), .B2(n16), .ZN(to_7[7])
         );
  LVT_AOI22HSV4 U106 ( .A1(ti_7[1]), .A2(ctro), .B1(t_i_2_out[1]), .B2(n16), 
        .ZN(n35) );
  LVT_CLKAND2HSV4 U107 ( .A1(t_i_2_out[15]), .A2(n16), .Z(n48) );
  LVT_NAND2HSV0 U108 ( .A1(ti_7[5]), .A2(ctro), .ZN(n36) );
  LVT_AOI22HSV4 U109 ( .A1(ti_7[16]), .A2(ctro), .B1(t_i_2_out[16]), .B2(n16), 
        .ZN(n39) );
  LVT_NAND2HSV12 U110 ( .A1(n101), .A2(l_t_i_1_in_0), .ZN(n89) );
  LVT_CLKAND2HSV4 U111 ( .A1(t_i_2_out[12]), .A2(n16), .Z(n55) );
  LVT_AO22HSV1 U112 ( .A1(mux_bq[28]), .A2(n33), .B1(b_out[28]), .B2(n90), .Z(
        mux_b[28]) );
  LVT_AO22HSV1 U113 ( .A1(mux_bq[29]), .A2(n33), .B1(b_out[29]), .B2(n90), .Z(
        mux_b[29]) );
  LVT_AO22HSV1 U114 ( .A1(mux_bq[30]), .A2(n33), .B1(b_out[30]), .B2(n90), .Z(
        mux_b[30]) );
  LVT_AO22HSV1 U115 ( .A1(n29), .A2(n33), .B1(b_out[31]), .B2(n90), .Z(
        mux_b[31]) );
  LVT_AOI22HSV4 U116 ( .A1(ti_7[13]), .A2(ctro), .B1(t_i_2_out[13]), .B2(n16), 
        .ZN(n40) );
  LVT_AOI22HSV4 U117 ( .A1(ti_7[9]), .A2(ctro), .B1(t_i_2_out[9]), .B2(n16), 
        .ZN(n41) );
  LVT_AOI22HSV4 U118 ( .A1(ti_7[29]), .A2(ctro), .B1(t_i_2_out[29]), .B2(n16), 
        .ZN(n42) );
  LVT_INHSV0SR U119 ( .I(n105), .ZN(n43) );
  LVT_INHSV2 U120 ( .I(n43), .ZN(t_i_2_out[7]) );
  LVT_INHSV0SR U121 ( .I(to_7[4]), .ZN(n45) );
  LVT_INHSV2 U122 ( .I(n45), .ZN(n46) );
  LVT_AO22HSV4 U123 ( .A1(ti_7[25]), .A2(ctro), .B1(t_i_2_out[25]), .B2(n16), 
        .Z(to_7[25]) );
  LVT_AND2HSV0RD U124 ( .A1(ti_7[15]), .A2(ctro), .Z(n47) );
  LVT_INHSV0SR U125 ( .I(l_t_i_1_in_0), .ZN(n102) );
  LVT_AND2HSV0RD U126 ( .A1(ti_7[19]), .A2(ctro), .Z(n50) );
  LVT_NAND2HSV0 U127 ( .A1(ti_7[8]), .A2(ctro), .ZN(n52) );
  LVT_AND2HSV0RD U128 ( .A1(ti_7[12]), .A2(ctro), .Z(n54) );
  LVT_AND2HSV0RD U129 ( .A1(ti_7[27]), .A2(ctro), .Z(n56) );
  LVT_AOI22HSV4 U130 ( .A1(ti_7[28]), .A2(ctro), .B1(t_i_2_out[28]), .B2(n16), 
        .ZN(n58) );
  LVT_AOI22HSV4 U131 ( .A1(ti_7[3]), .A2(ctro), .B1(t_i_2_out[3]), .B2(n16), 
        .ZN(n59) );
  LVT_AOI22HSV4 U132 ( .A1(ti_7[2]), .A2(ctro), .B1(t_i_2_out[2]), .B2(n16), 
        .ZN(n60) );
  LVT_AOI22HSV4 U133 ( .A1(ti_7[11]), .A2(ctro), .B1(t_i_2_out[11]), .B2(n16), 
        .ZN(n61) );
  LVT_AOI22HSV4 U134 ( .A1(ti_7[0]), .A2(ctro), .B1(t_i_2_out[0]), .B2(n16), 
        .ZN(n62) );
  LVT_NAND2HSV0 U135 ( .A1(ti_7[4]), .A2(ctro), .ZN(n64) );
  LVT_AND2HSV0RD U136 ( .A1(ti_7[18]), .A2(ctro), .Z(n66) );
  LVT_NAND2HSV0 U137 ( .A1(ti_7[26]), .A2(ctro), .ZN(n68) );
  LVT_NAND2HSV0 U138 ( .A1(ti_7[6]), .A2(ctro), .ZN(n70) );
  LVT_BUFHSV2RT U139 ( .I(n33), .Z(n83) );
  LVT_NAND2HSV0 U140 ( .A1(ti_7[14]), .A2(ctro), .ZN(n84) );
  LVT_INHSV0SR U141 ( .I(n104), .ZN(n86) );
  LVT_INHSV2 U142 ( .I(n86), .ZN(t_i_2_out[17]) );
  LVT_AO22HSV4 U143 ( .A1(ti_7[21]), .A2(ctro), .B1(t_i_2_out[21]), .B2(n16), 
        .Z(to_7[21]) );
  LVT_AO22HSV4 U144 ( .A1(ti_7[30]), .A2(ctro), .B1(t_i_2_out[30]), .B2(n15), 
        .Z(to_7[30]) );
endmodule


module regist_32bit_5 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3, n4;

  LVT_DRNQHSV4 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV4 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV4 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV4 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n3), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n3), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n3), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n3), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n3), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n3), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n3), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n3), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_INHSV2 U3 ( .I(n4), .ZN(n2) );
  LVT_INHSV2 U4 ( .I(n4), .ZN(n1) );
  LVT_INHSV2 U5 ( .I(rstn), .ZN(n4) );
  LVT_INHSV2 U6 ( .I(n4), .ZN(n3) );
endmodule


module regist_32bit_4 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV2 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n2), .Q(out[31]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n2), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n2), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n2), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n2), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n2), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n1), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n1), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n1), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n1), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n1), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n1), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n1), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n2), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n2), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n2), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n2), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_32bit_3 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3, n4;

  LVT_DRNQHSV4 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV4 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV4 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV4 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV4 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV4 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV4 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n3), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n3), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n3), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n3), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n3), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n3), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n3), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n3), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_INHSV2 U3 ( .I(n4), .ZN(n2) );
  LVT_INHSV2 U4 ( .I(n4), .ZN(n1) );
  LVT_INHSV2 U5 ( .I(rstn), .ZN(n4) );
  LVT_INHSV2 U6 ( .I(n4), .ZN(n3) );
endmodule


module regist_1bit_3 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_1bit_2 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_31bit_3 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n1), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n1), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n2), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n2), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n2), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n2), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n2), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n2), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n1), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n1), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n1), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n1), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n1), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n1), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n1), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n2), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n2), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n2), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_INHSV2 U3 ( .I(n3), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n2) );
endmodule


module regist_31bit_2 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n1), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n2), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(rstn), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n1), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n2), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n1), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n1), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n2), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n2), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n2), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n2), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(rstn), .Q(out[11])
         );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n2), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n2), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n1), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n1), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n1), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n2), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n2), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_INHSV2 U3 ( .I(n3), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n2) );
endmodule


module regist_1bit_1 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV4 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_32bit_2 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3, n4;

  LVT_DRNQHSV4 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n3), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n3), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n1), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n1), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n1), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n3), .Q(out[0]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n2), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n2), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n2), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n2), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n2), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n2), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n2), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n2), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n3), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n3), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n3), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n3), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n3), .Q(out[15]) );
  LVT_INHSV2 U3 ( .I(n4), .ZN(n2) );
  LVT_INHSV2 U4 ( .I(rstn), .ZN(n4) );
  LVT_INHSV2 U5 ( .I(n4), .ZN(n3) );
  LVT_INHSV2 U6 ( .I(n4), .ZN(n1) );
endmodule


module regist_1bit_0 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV2 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module regist_31bit_1 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2;

  LVT_DRNQHSV1 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(rstn), .Q(out[0]) );
  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(rstn), .Q(out[30])
         );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(rstn), .Q(out[26])
         );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(rstn), .Q(out[24])
         );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n1), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n1), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(rstn), .Q(out[10])
         );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(rstn), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(rstn), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(rstn), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(rstn), .Q(out[11])
         );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n1), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n1), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n1), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(rstn), .Q(out[1]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(rstn), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(rstn), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n1), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(rstn), .Q(out[2]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(rstn), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n1), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n1), .Q(out[12]) );
  LVT_INHSV0SR U3 ( .I(rstn), .ZN(n2) );
  LVT_INHSV2 U4 ( .I(n2), .ZN(n1) );
endmodule


module cell_3_961 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_4_30 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_29 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_28 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_27 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_26 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_25 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_24 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_23 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_22 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_21 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_20 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_19 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_18 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_17 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_16 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_15 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_14 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR3HSV1 U1 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
endmodule


module cell_4_13 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
endmodule


module cell_4_12 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV2 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(n7) );
endmodule


module cell_4_11 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_10 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_9 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_8 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_4_7 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_4_6 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_4_5 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n2) );
  LVT_XOR3HSV1 U2 ( .A1(n5), .A2(n4), .A3(n2), .Z(t_i_out) );
endmodule


module cell_4_4 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XOR2HSV0 U3 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_4_3 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_NAND2HSV0 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_4_2 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n8) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(n7) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_4_1 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n1, n5, n6, n7, n8, n9;

  LVT_OAI21HSV2 U1 ( .A1(n1), .A2(n7), .B(n5), .ZN(n9) );
  LVT_NAND2HSV0P5 U2 ( .A1(n7), .A2(n1), .ZN(n5) );
  LVT_INHSV0SR U3 ( .I(n8), .ZN(n1) );
  LVT_NAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XNOR2HSV1 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n7) );
  LVT_XNOR2HSV4 U7 ( .A1(n6), .A2(n9), .ZN(t_i_out) );
endmodule


module cell_4_0 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in;
  output t_i_out;
  wire   n2, n3, n5, n6;

  LVT_XOR2HSV0 U5 ( .A1(t_i_2_in), .A2(t_i_1_in), .Z(n6) );
  LVT_XOR2HSV4 U1 ( .A1(n5), .A2(n2), .Z(n3) );
  LVT_CLKNAND2HSV4 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_CLKAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .Z(n2) );
  LVT_XNOR2HSV4 U4 ( .A1(n6), .A2(n3), .ZN(t_i_out) );
endmodule


module row_1_0 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_2_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [31:0] t_i_1_in;
  input [30:0] t_i_2_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_3_961 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[0]) );
  cell_4_30 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[1]), .t_i_2_in(t_i_2_in[0]), .t_i_out(t_i_1_out[1])
         );
  cell_4_29 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[2]), .t_i_2_in(t_i_2_in[1]), .t_i_out(t_i_1_out[2])
         );
  cell_4_28 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_2_in(t_i_2_in[2]), .t_i_out(t_i_1_out[3])
         );
  cell_4_27 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_2_in(t_i_2_in[3]), .t_i_out(t_i_1_out[4])
         );
  cell_4_26 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_2_in(t_i_2_in[4]), .t_i_out(t_i_1_out[5])
         );
  cell_4_25 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_2_in(t_i_2_in[5]), .t_i_out(t_i_1_out[6])
         );
  cell_4_24 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_2_in(t_i_2_in[6]), .t_i_out(t_i_1_out[7])
         );
  cell_4_23 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_2_in(t_i_2_in[7]), .t_i_out(t_i_1_out[8])
         );
  cell_4_22 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[9]), .t_i_2_in(t_i_2_in[8]), .t_i_out(t_i_1_out[9])
         );
  cell_4_21 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[10]), .t_i_2_in(t_i_2_in[9]), .t_i_out(
        t_i_1_out[10]) );
  cell_4_20 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[11]), .t_i_2_in(t_i_2_in[10]), .t_i_out(
        t_i_1_out[11]) );
  cell_4_19 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[12]), .t_i_2_in(t_i_2_in[11]), .t_i_out(
        t_i_1_out[12]) );
  cell_4_18 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[13]), .t_i_2_in(t_i_2_in[12]), .t_i_out(
        t_i_1_out[13]) );
  cell_4_17 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[14]), .t_i_2_in(t_i_2_in[13]), .t_i_out(
        t_i_1_out[14]) );
  cell_4_16 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[15]), .t_i_2_in(t_i_2_in[14]), .t_i_out(
        t_i_1_out[15]) );
  cell_4_15 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[16]), .t_i_2_in(t_i_2_in[15]), .t_i_out(
        t_i_1_out[16]) );
  cell_4_14 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[17]), .t_i_2_in(t_i_2_in[16]), .t_i_out(
        t_i_1_out[17]) );
  cell_4_13 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[18]), .t_i_2_in(t_i_2_in[17]), .t_i_out(
        t_i_1_out[18]) );
  cell_4_12 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[19]), .t_i_2_in(t_i_2_in[18]), .t_i_out(
        t_i_1_out[19]) );
  cell_4_11 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_2_in(t_i_2_in[19]), .t_i_out(
        t_i_1_out[20]) );
  cell_4_10 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_2_in(t_i_2_in[20]), .t_i_out(
        t_i_1_out[21]) );
  cell_4_9 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_2_in(t_i_2_in[21]), .t_i_out(
        t_i_1_out[22]) );
  cell_4_8 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_2_in(t_i_2_in[22]), .t_i_out(
        t_i_1_out[23]) );
  cell_4_7 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_2_in(t_i_2_in[23]), .t_i_out(
        t_i_1_out[24]) );
  cell_4_6 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_2_in(t_i_2_in[24]), .t_i_out(
        t_i_1_out[25]) );
  cell_4_5 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_2_in(t_i_2_in[25]), .t_i_out(
        t_i_1_out[26]) );
  cell_4_4 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_2_in(t_i_2_in[26]), .t_i_out(
        t_i_1_out[27]) );
  cell_4_3 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_2_in(t_i_2_in[27]), .t_i_out(
        t_i_1_out[28]) );
  cell_4_2 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_2_in(t_i_2_in[28]), .t_i_out(
        t_i_1_out[29]) );
  cell_4_1 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_2_in(t_i_2_in[29]), .t_i_out(
        t_i_1_out[30]) );
  cell_4_0 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[31]), .t_i_2_in(t_i_2_in[30]), .t_i_out(
        t_i_2_out) );
  LVT_INHSV0P5SR U1 ( .I(t_m_1_in), .ZN(n2) );
  LVT_INHSV2 U2 ( .I(n2), .ZN(n3) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n1) );
  LVT_BUFHSV2RQ U4 ( .I(n1), .Z(n4) );
endmodule


module cell_2_30 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_960 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_959 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_958 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_957 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_956 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_955 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_954 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_953 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_952 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_951 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_950 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_949 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_948 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_947 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_946 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_945 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_944 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_943 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_942 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_941 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_940 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_939 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_938 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_937 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_936 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_935 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_934 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_933 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_932 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_931 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4, n5, n6, n7, n8;

  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_CLKAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .Z(n6) );
  LVT_NAND2HSV2 U4 ( .A1(n2), .A2(n3), .ZN(n5) );
  LVT_NAND2HSV0 U5 ( .A1(n8), .A2(n7), .ZN(n4) );
  LVT_NAND2HSV2 U6 ( .A1(n4), .A2(n5), .ZN(t_i_out) );
  LVT_CLKNHSV0P5 U7 ( .I(n8), .ZN(n2) );
  LVT_INHSV2 U8 ( .I(n7), .ZN(n3) );
endmodule


module cell_3_930 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;

  LVT_CLKNAND2HSV3 U1 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNAND2HSV8 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n13) );
  LVT_INHSV2 U3 ( .I(n11), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(n9), .A2(n10), .ZN(n11) );
  LVT_INHSV2 U5 ( .I(n13), .ZN(n2) );
  LVT_INHSV2 U6 ( .I(t_i_1_in), .ZN(n8) );
  LVT_NAND2HSV2 U7 ( .A1(n12), .A2(n8), .ZN(n9) );
  LVT_NAND2HSV1 U8 ( .A1(n7), .A2(t_i_1_in), .ZN(n10) );
  LVT_NAND2HSV2 U9 ( .A1(n13), .A2(n4), .ZN(n5) );
  LVT_CLKNAND2HSV3 U10 ( .A1(n2), .A2(n11), .ZN(n6) );
  LVT_CLKNHSV0 U11 ( .I(n12), .ZN(n7) );
  LVT_NAND2HSV0 U12 ( .A1(b_in), .A2(a_in), .ZN(n12) );
endmodule


module row_other_30 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_30 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_960 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_959 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_958 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_957 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_956 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_955 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_954 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_953 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_952 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_951 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_950 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_949 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_948 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_947 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_946 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_945 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_944 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_943 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_942 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_941 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_940 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_939 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_938 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_937 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_936 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_935 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_934 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_933 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_932 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_931 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_930 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV6 U1 ( .I(n1), .ZN(n2) );
  LVT_CLKNHSV2 U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_29 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_929 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_928 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_927 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_926 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_925 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_924 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_923 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_922 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_921 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_920 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_919 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_918 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_917 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_916 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_915 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_914 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_913 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_912 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_911 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_910 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_909 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_908 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_907 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_906 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_905 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n5), .A2(n6), .Z(t_i_out) );
endmodule


module cell_3_904 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_903 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_902 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_901 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_900 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_899 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(n5), .A2(n6), .ZN(n9) );
  LVT_NAND2HSV4 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_CLKXOR2HSV4 U4 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U5 ( .A1(n7), .A2(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV2 U6 ( .A1(n8), .A2(n4), .ZN(n6) );
  LVT_CLKNHSV1 U7 ( .I(t_i_1_in), .ZN(n4) );
  LVT_INHSV2 U8 ( .I(n8), .ZN(n7) );
endmodule


module row_other_29 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_29 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_929 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_928 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_927 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_926 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_925 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_924 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_923 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_922 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_921 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_920 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_919 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_918 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_917 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_916 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_915 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_914 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_913 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_912 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_911 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_910 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_909 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_908 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_907 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_906 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_905 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_904 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_903 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_902 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_901 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_900 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_899 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_28 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_898 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_897 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_896 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_895 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_894 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_893 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_892 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_891 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_890 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_889 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_888 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_887 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_886 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_885 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_884 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_883 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_882 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_881 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_880 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_879 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_878 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_877 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_876 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_875 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_874 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_873 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_872 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_871 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_870 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_869 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV4 U1 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV0P5 U4 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U6 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0SR U7 ( .I(n8), .ZN(n4) );
  LVT_INHSV2 U8 ( .I(t_i_1_in), .ZN(n5) );
endmodule


module cell_3_868 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_OAI21HSV2 U1 ( .A1(n6), .A2(n4), .B(n2), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKNAND2HSV1 U4 ( .A1(n6), .A2(n4), .ZN(n2) );
  LVT_XNOR2HSV4 U5 ( .A1(n5), .A2(t_i_1_in), .ZN(n4) );
endmodule


module row_other_28 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1;

  cell_2_28 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_898 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_897 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_896 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_895 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_894 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_893 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_892 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_891 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_890 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_889 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_888 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_887 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_886 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_885 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_884 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_883 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_882 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_881 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_880 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_879 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_878 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_877 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_876 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_875 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_874 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_873 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_872 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_871 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_870 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_869 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_868 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV2RT U1 ( .I(t_m_1_in), .Z(n1) );
endmodule


module cell_2_27 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_867 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_866 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_865 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_864 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_863 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_862 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_861 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_860 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_859 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_858 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_857 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_856 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_855 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_854 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_853 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_852 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_851 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_850 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_849 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_848 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_847 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_846 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV0P5 U1 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U5 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0SR U6 ( .I(n8), .ZN(n4) );
  LVT_CLKNHSV0P5 U7 ( .I(t_i_1_in), .ZN(n5) );
  LVT_XOR2HSV2 U8 ( .A1(n10), .A2(n9), .Z(t_i_out) );
endmodule


module cell_3_845 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_844 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_843 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_842 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_841 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_840 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_839 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_838 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_837 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_27 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_27 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_867 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_866 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_865 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_864 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_863 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_862 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_861 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_860 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_859 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_858 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_857 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_856 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_855 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_854 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_853 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_852 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_851 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_850 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_849 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_848 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_847 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_846 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_845 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_844 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_843 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_842 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_841 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_840 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_839 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_838 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_837 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV6 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV2 U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_26 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_836 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_835 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_834 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_833 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_832 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_831 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_830 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_829 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_828 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_827 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_826 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_825 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_824 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_823 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_822 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_821 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_820 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_819 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_818 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_817 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_816 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_815 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_814 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_813 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_812 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_811 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV3 U1 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0P5 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
  LVT_INHSV0SR U5 ( .I(n10), .ZN(n4) );
  LVT_INHSV2P5 U6 ( .I(n9), .ZN(n5) );
  LVT_NAND2HSV0 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_XOR2HSV2 U8 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
endmodule


module cell_3_810 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_809 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_808 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_807 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_806 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_26 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_26 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_836 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_835 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_834 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_833 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_832 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_831 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_830 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_829 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_828 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_827 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_826 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_825 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_824 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_823 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_822 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_821 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_820 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_819 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_818 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_817 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_816 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_815 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_814 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_813 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_812 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_811 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_810 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_809 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_808 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_807 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_806 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV2RT U1 ( .I(n3), .Z(n1) );
  LVT_INHSV4SR U2 ( .I(n2), .ZN(n3) );
  LVT_INHSV0SR U3 ( .I(t_m_1_in), .ZN(n2) );
endmodule


module cell_2_25 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_805 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_804 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_803 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_802 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_801 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_800 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_799 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_798 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_797 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_796 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_795 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_794 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_793 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_792 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_791 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_790 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_789 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_788 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_787 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_786 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_785 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_784 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_783 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_782 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV1 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_NAND2HSV0 U4 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_INHSV0SR U5 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_781 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(t_i_1_in), .Z(n7) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV1 U1 ( .A1(n4), .A2(n7), .B(n5), .ZN(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(n4), .A2(n7), .ZN(n5) );
  LVT_INHSV0SR U5 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_780 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_779 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV1 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV0P5 U5 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_778 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_777 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV1 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_776 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV4 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_775 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module row_other_25 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_2_25 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_805 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_804 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_803 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_802 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_801 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_800 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_799 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_798 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_797 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_796 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_795 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_794 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_793 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_792 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_791 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_790 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_789 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_788 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_787 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_786 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_785 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_784 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_783 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_782 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_781 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_780 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_779 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_778 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_777 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_776 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_775 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV4 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV2 U2 ( .I(n4), .ZN(n3) );
  LVT_INHSV0SR U3 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV0SR U4 ( .I(n2), .ZN(n4) );
endmodule


module cell_2_24 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_774 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_773 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_772 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_771 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_770 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_769 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_768 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_767 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_766 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_765 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_764 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_763 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_762 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_761 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_760 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_759 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_758 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_757 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_756 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_755 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_754 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_753 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_752 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_751 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_750 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_749 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_748 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U3 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV2 U5 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_747 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_746 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_745 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_744 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_24 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_24 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_774 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_773 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_772 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_771 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_770 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_769 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_768 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_767 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_766 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_765 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_764 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_763 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_762 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_761 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_760 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_759 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_758 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_757 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_756 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_755 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_754 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_753 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_752 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_751 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_750 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_749 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_748 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_747 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_746 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_745 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_744 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV4 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV2 U2 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2SR U3 ( .I(n1), .ZN(n3) );
endmodule


module cell_2_23 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_743 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_742 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_741 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_740 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_739 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_738 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_737 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_736 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_735 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_734 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_733 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_732 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_731 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_730 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_729 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_728 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_727 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_726 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_725 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_724 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_723 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_722 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_721 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_720 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_719 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_718 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_717 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_716 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(t_i_1_in), .A2(n4), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_715 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_CLKNAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV2 U5 ( .I(n6), .ZN(n4) );
  LVT_XOR2HSV2 U6 ( .A1(n7), .A2(n8), .Z(t_i_out) );
endmodule


module cell_3_714 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_713 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module row_other_23 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_23 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_743 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_742 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_741 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_740 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_739 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_738 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_737 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_736 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_735 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_734 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_733 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_732 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_731 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_730 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_729 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_728 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_727 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_726 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_725 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_724 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_723 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_722 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_721 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_720 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_719 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_718 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_717 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_716 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_715 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_714 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_713 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV0 U1 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U2 ( .I(t_m_1_in), .ZN(n2) );
  LVT_CLKNHSV6 U3 ( .I(n2), .ZN(n3) );
endmodule


module cell_2_22 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_712 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_711 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_710 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_709 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_708 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_707 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_706 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_705 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_704 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_703 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_702 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_701 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_700 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_699 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_698 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_697 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_696 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_695 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_694 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_693 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_692 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_691 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_690 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_689 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_688 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_687 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_686 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_685 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_684 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV2 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
endmodule


module cell_3_683 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_682 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_NAND2HSV0P5 U1 ( .A1(n6), .A2(n4), .ZN(n2) );
  LVT_OAI21HSV2 U2 ( .A1(n6), .A2(n4), .B(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XNOR2HSV4 U5 ( .A1(n5), .A2(t_i_1_in), .ZN(n4) );
endmodule


module row_other_22 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_22 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_712 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_711 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_710 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_709 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_708 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_707 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_706 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_705 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_704 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_703 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_702 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_701 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_700 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_699 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_698 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_697 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_696 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_695 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_694 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_693 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_692 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_691 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_690 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_689 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_688 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_687 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_686 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_685 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_684 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_683 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_682 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV6 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV2 U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_21 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_681 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_680 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_679 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_678 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_677 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_676 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_675 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_674 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_673 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_672 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_671 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_670 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_669 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_668 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_667 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_666 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_665 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_664 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_663 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_662 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_661 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_660 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_659 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_658 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_657 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_656 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_655 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_NAND2HSV2 U1 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U2 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0 U3 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_CLKNHSV0 U5 ( .I(n8), .ZN(n4) );
  LVT_CLKNHSV2 U6 ( .I(t_i_1_in), .ZN(n5) );
  LVT_XOR2HSV0 U7 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV0 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_654 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_653 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_652 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_OAI21HSV2 U1 ( .A1(n6), .A2(n4), .B(n2), .ZN(t_i_out) );
  LVT_NAND2HSV0 U2 ( .A1(n6), .A2(n4), .ZN(n2) );
  LVT_XNOR2HSV4 U4 ( .A1(n5), .A2(t_i_1_in), .ZN(n4) );
  LVT_NAND2HSV0 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_651 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_21 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_21 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_681 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_680 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_679 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_678 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_677 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_676 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_675 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_674 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_673 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_672 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_671 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_670 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_669 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_668 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_667 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_666 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_665 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_664 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_663 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_662 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_661 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_660 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_659 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_658 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_657 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_656 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_655 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_654 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_653 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_652 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_651 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2SR U1 ( .I(n2), .ZN(n1) );
  LVT_INHSV0SR U2 ( .I(t_m_1_in), .ZN(n2) );
endmodule


module cell_2_20 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_650 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_649 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_648 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_647 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_646 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_645 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_644 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_643 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_642 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_641 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_640 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_639 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_638 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_637 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_636 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_635 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_634 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_633 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_632 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_631 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_630 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_629 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_628 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_627 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_626 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_625 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_624 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_623 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_622 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_621 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_620 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_20 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_20 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_650 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_649 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_648 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_647 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_646 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_645 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_644 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_643 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_642 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_641 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_640 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_639 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_638 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_637 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_636 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_635 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_634 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_633 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_632 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_631 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_630 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_629 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_628 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_627 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_626 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_625 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_624 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_623 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_622 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_621 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_620 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_19 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_619 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_618 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_617 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_616 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_615 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_614 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_613 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_612 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_611 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_610 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_609 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_608 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_607 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_606 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_605 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_604 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_603 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_602 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_601 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_600 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_599 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_598 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_597 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_596 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_595 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_594 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_593 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_592 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_591 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_590 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_589 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV4 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module row_other_19 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_19 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_619 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_618 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_617 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_616 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_615 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_614 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_613 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_612 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_611 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_610 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_609 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_608 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_607 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_606 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_605 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_604 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_603 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_602 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_601 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_600 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_599 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_598 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_597 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_596 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_595 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_594 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_593 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_592 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_591 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_590 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_589 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV4 U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV10 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_18 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_588 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_587 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_586 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_585 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_584 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_583 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_582 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_581 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_580 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_579 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_578 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_577 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_576 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_575 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_574 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_573 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_572 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_571 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_570 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_569 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_568 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_567 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_566 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_565 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_564 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_563 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_562 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_561 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_560 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_559 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV4 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_CLKXOR2HSV4 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_558 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_18 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1;

  cell_2_18 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_588 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_587 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_586 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_585 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_584 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_583 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_582 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_581 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_580 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_579 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_578 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_577 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_576 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_575 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_574 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_573 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_572 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_571 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_570 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_569 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_568 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_567 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_566 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_565 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_564 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_563 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_562 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_561 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_560 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_559 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_558 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV6 U1 ( .I(t_m_1_in), .Z(n1) );
endmodule


module cell_2_17 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_557 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_556 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_555 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_554 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_553 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_552 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_551 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_550 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_549 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_548 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_547 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_546 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_545 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_544 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_543 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_542 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_541 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_540 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_539 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_538 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_537 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_536 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_535 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_534 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_533 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_532 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_531 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_530 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_529 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_528 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_527 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV4 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV4 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module row_other_17 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_17 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_557 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_556 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_555 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_554 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_553 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_552 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_551 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_550 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_549 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_548 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_547 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_546 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_545 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_544 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_543 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_542 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_541 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_540 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_539 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_538 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_537 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_536 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_535 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_534 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_533 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_532 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_531 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_530 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_529 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_528 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_527 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV8 U1 ( .I(n1), .ZN(n2) );
  LVT_CLKNHSV4 U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_16 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_526 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_525 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_524 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_523 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_522 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_521 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_520 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_519 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_518 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_517 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_516 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_515 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_514 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_513 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_512 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_511 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_510 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_509 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_508 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_507 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_506 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_505 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_504 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_503 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_502 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_501 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_500 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_499 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_498 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_497 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_496 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_16 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_16 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_526 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_525 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_524 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_523 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_522 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_521 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_520 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_519 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_518 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_517 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_516 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_515 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_514 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_513 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_512 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_511 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_510 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_509 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_508 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_507 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_506 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_505 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_504 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_503 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_502 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_501 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_500 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_499 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_498 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_497 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_496 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_15 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_495 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_494 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_493 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_492 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_491 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_490 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_489 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_488 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_487 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_486 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_485 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_484 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_483 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_482 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_481 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_480 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_479 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_478 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_477 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_476 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_475 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_474 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_473 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_472 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_471 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_470 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_469 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_468 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_467 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_466 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_465 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n3, n4;

  LVT_CLKAND2HSV2 U1 ( .A1(b_in), .A2(a_in), .Z(n2) );
  LVT_XOR2HSV4 U2 ( .A1(n2), .A2(t_i_1_in), .Z(n3) );
  LVT_CLKNAND2HSV3 U3 ( .A1(t_m_1_in), .A2(g_in), .ZN(n4) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(n3), .ZN(t_i_out) );
endmodule


module row_other_15 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_15 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_495 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_494 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_493 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_492 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_491 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_490 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_489 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_488 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_487 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_486 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_485 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_484 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_483 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_482 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_481 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_480 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_479 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_478 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_477 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_476 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_475 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_474 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_473 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_472 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_471 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_470 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_469 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_468 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_467 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_466 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_465 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV10 U1 ( .I(n2), .ZN(n1) );
  LVT_INHSV4SR U2 ( .I(t_m_1_in), .ZN(n2) );
endmodule


module cell_2_14 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_464 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_463 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_462 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_461 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_460 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_459 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_458 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_457 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_456 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_455 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_454 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_453 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_452 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_451 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_450 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_449 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_448 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_447 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_446 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_445 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_444 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_443 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_442 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_441 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_440 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_439 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_438 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_437 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_436 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_435 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNHSV0P5 U1 ( .I(n9), .ZN(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n8), .A2(t_i_1_in), .Z(n9) );
  LVT_INHSV2 U4 ( .I(n10), .ZN(n4) );
  LVT_NAND2HSV2 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_NAND2HSV0P5 U6 ( .A1(n10), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U7 ( .A1(n4), .A2(n9), .ZN(n7) );
  LVT_NAND2HSV2 U8 ( .A1(n6), .A2(n7), .ZN(t_i_out) );
endmodule


module cell_3_434 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV8 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_14 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_14 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_464 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_463 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_462 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_461 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_460 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_459 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_458 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_457 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_456 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_455 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_454 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_453 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_452 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_451 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_450 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_449 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_448 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_447 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_446 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_445 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_444 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_443 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_442 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_441 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_440 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_439 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_438 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_437 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_436 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_435 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_434 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_13 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_433 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_432 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_431 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_430 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_429 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_428 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_427 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_426 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_425 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_424 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_423 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_422 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_421 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_420 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_419 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_418 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_417 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_416 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_415 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_414 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_413 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_412 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_411 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_410 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_409 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_408 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_407 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_406 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_405 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module cell_3_404 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV4 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_403 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV2 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNHSV2 U4 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV3 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV0P5 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV3SR U7 ( .I(n9), .ZN(n2) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_13 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_13 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_433 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_432 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_431 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_430 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_429 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_428 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_427 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_426 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_425 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_424 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_423 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_422 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_421 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_420 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_419 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_418 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_417 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_416 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_415 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_414 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_413 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_412 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_411 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_410 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_409 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_408 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_407 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_406 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_405 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_404 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_403 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV1 U1 ( .I(t_m_1_in), .ZN(n1) );
  LVT_CLKNHSV4 U2 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_12 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_402 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_401 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_400 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_399 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_398 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_397 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_396 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_395 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_394 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_393 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_392 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_391 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_390 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_389 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_388 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_387 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_386 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_385 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_384 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_383 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_382 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_381 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_380 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_379 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_378 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_377 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_376 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_375 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_374 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_373 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_372 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_NAND2HSV2 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2 U4 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV0P5 U5 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV2 U6 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV2 U7 ( .I(n9), .ZN(n2) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_12 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_12 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_402 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_401 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_400 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_399 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_398 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_397 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_396 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_395 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_394 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_393 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_392 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_391 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_390 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_389 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_388 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_387 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_386 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_385 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_384 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_383 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_382 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_381 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_380 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_379 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_378 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_377 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_376 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_375 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_374 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_373 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_372 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV1SR U1 ( .I(t_m_1_in), .ZN(n2) );
  LVT_CLKNHSV8 U2 ( .I(n2), .ZN(n1) );
endmodule


module cell_2_11 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_371 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_370 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_369 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_368 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_367 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_366 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_365 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_364 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_363 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_362 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_361 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_360 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_359 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_358 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_357 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_356 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_355 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_354 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_353 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_352 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_351 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_350 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_349 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_348 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_347 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_346 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_345 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_344 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_343 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_342 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_341 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_11 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_11 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_371 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_370 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_369 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_368 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_367 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_366 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_365 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_364 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_363 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_362 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_361 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_360 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_359 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_358 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_357 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_356 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_355 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_354 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_353 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_352 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_351 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_350 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_349 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_348 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_347 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_346 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_345 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_344 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_343 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_342 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_341 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_10 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_340 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_339 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_338 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_337 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_336 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_335 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_334 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_333 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_332 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_331 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_330 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_329 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_328 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_327 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_326 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_325 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_324 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_323 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_322 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_321 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_320 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_319 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_318 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_317 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_316 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_315 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_314 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_313 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_312 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV1 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U5 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_311 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_310 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n7) );
  LVT_NAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_IOA21HSV2 U2 ( .A1(n8), .A2(n6), .B(n5), .ZN(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(n2), .A2(n4), .ZN(n5) );
  LVT_XNOR2HSV1 U5 ( .A1(n7), .A2(t_i_1_in), .ZN(n6) );
  LVT_INHSV2SR U6 ( .I(n8), .ZN(n2) );
  LVT_INHSV2SR U7 ( .I(n6), .ZN(n4) );
endmodule


module row_other_10 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_10 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_340 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_339 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_338 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_337 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_336 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_335 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_334 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n3), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_333 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_332 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_331 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_330 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_329 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_328 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_327 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_326 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_325 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_324 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_323 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_322 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_321 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_320 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n3), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_319 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_318 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_317 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_316 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_315 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_314 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_313 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_312 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_311 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_310 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV0P5 U1 ( .I(t_m_1_in), .ZN(n2) );
  LVT_INHSV2 U2 ( .I(n2), .ZN(n1) );
  LVT_INHSV2 U3 ( .I(n2), .ZN(n3) );
endmodule


module cell_2_9 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_309 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_308 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_307 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_306 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_305 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_304 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_303 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_302 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_301 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_300 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_299 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_298 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_297 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_296 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_295 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_294 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_293 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_292 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_291 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_290 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_289 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_288 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_287 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_286 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_285 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_284 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_XOR2HSV0 U4 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_283 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_282 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_281 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_280 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_279 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n4), .ZN(n2) );
endmodule


module row_other_9 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_9 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_309 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_308 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_307 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_306 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_305 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_304 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_303 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_302 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_301 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_300 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_299 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_298 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_297 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_296 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_295 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_294 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_293 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_292 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_291 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_290 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_289 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_288 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_287 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_286 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_285 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_284 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_283 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_282 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_281 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_280 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_279 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV12 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV6SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_8 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_278 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_277 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_276 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_275 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_274 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_273 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_272 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_271 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_270 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_269 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_268 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_267 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_266 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_265 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_264 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_263 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_262 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_261 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_260 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_259 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_258 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_257 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_256 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_255 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_254 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_253 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_252 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_251 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_250 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_249 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKXOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_248 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_8 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_8 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_278 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_277 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_276 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_275 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_274 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_273 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_272 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_271 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_270 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_269 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_268 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_267 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_266 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_265 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_264 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_263 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_262 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_261 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_260 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_259 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_258 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_257 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_256 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_255 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_254 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_253 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_252 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_251 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_250 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_249 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_248 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV4 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV2 U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_7 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_247 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_246 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_245 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_244 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_243 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_242 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_241 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_240 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_239 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_238 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_237 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_236 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_235 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_234 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_233 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_232 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_231 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_230 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_229 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_228 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_227 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_226 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_225 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_224 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_223 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_222 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_221 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_220 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV2 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_219 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
  LVT_XOR2HSV0 U2 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV2 U4 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U6 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV2 U7 ( .I(n8), .ZN(n4) );
  LVT_INHSV2 U8 ( .I(t_i_1_in), .ZN(n5) );
endmodule


module cell_3_218 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_OAI21HSV1 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_NAND2HSV0P5 U3 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U4 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV2 U5 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_XOR2HSV2 U6 ( .A1(n8), .A2(n7), .Z(t_i_out) );
endmodule


module cell_3_217 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_INHSV2SR U2 ( .I(n9), .ZN(n2) );
  LVT_XNOR2HSV4 U4 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV1 U6 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV2 U7 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV2 U8 ( .I(n7), .ZN(n4) );
endmodule


module row_other_7 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3;

  cell_2_7 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_247 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_246 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_245 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_244 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_243 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_242 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_241 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_240 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_239 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_238 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_237 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_236 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_235 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_234 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_233 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_232 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_231 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_230 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_229 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_228 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_227 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_226 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_225 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_224 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_223 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_222 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_221 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_220 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_219 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_218 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_217 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2SR U1 ( .I(t_m_1_in), .ZN(n3) );
  LVT_CLKNHSV4 U2 ( .I(n3), .ZN(n2) );
  LVT_INHSV1SR U3 ( .I(n3), .ZN(n1) );
endmodule


module cell_2_6 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_216 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_215 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_214 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_213 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_212 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_211 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_210 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_209 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_208 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_207 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_206 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_205 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_204 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_203 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_202 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_201 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_200 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_199 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_198 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_197 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_196 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_195 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_194 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_193 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_192 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_191 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_190 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_189 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_CLKNAND2HSV1 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_188 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_187 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV2 U3 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV0 U5 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(b_in), .A2(a_in), .ZN(n6) );
endmodule


module cell_3_186 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_6 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_6 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_216 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_215 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_214 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_213 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_212 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_211 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_210 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_209 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_208 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_207 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_206 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_205 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_204 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_203 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_202 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_201 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_200 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_199 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_198 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_197 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_196 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_195 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_194 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_193 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_192 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_191 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_190 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_189 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_188 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_187 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_186 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_5 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_185 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_184 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_183 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_182 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_181 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_180 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_179 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_178 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_177 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_176 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_175 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_174 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_173 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_172 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_171 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_170 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_169 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_168 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_167 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_166 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_165 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_164 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_163 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_162 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_161 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_160 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_159 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_158 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_157 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_156 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV2 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_155 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_NAND2HSV2 U1 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_INHSV2SR U2 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNHSV0P5 U5 ( .I(n9), .ZN(n2) );
  LVT_NAND2HSV2 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV4 U7 ( .A1(t_i_1_in), .A2(n8), .ZN(n7) );
  LVT_NAND2HSV0P5 U8 ( .A1(n9), .A2(n7), .ZN(n5) );
endmodule


module row_other_5 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_2_5 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_out(t_i_1_out[0]) );
  cell_3_185 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_184 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_183 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_182 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_181 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_180 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_179 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_178 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_177 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_176 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_175 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_174 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_173 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n4), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_172 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n4), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_171 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n4), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_170 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n4), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_169 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_168 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_167 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_166 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_165 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_164 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_163 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_162 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(n4), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_161 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(n1), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_160 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_159 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(n4), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_158 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_157 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_156 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_155 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV2P5 U1 ( .I(n3), .ZN(n4) );
  LVT_INHSV2 U2 ( .I(n3), .ZN(n1) );
  LVT_INHSV2 U3 ( .I(n3), .ZN(n2) );
  LVT_INHSV2SR U4 ( .I(t_m_1_in), .ZN(n3) );
endmodule


module cell_2_4 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_154 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_153 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_152 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_151 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_150 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_149 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_148 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_147 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_146 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_145 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_144 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_143 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_142 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_141 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_140 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_139 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_138 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_137 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_136 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_135 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_134 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_133 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_132 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_131 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_130 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_129 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_128 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_127 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_126 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_125 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNHSV2 U1 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV0P5 U2 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_CLKNAND2HSV3 U4 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_CLKNAND2HSV3 U5 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_CLKNHSV2 U6 ( .I(n9), .ZN(n2) );
  LVT_XNOR2HSV1 U7 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV0 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
endmodule


module cell_3_124 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV1 U1 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV2 U2 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_INHSV2P5 U5 ( .I(n9), .ZN(n2) );
  LVT_INHSV2 U6 ( .I(n7), .ZN(n4) );
  LVT_NAND2HSV2 U7 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_4 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2;

  cell_2_4 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_154 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_153 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_152 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_151 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_150 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_149 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_148 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_147 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_146 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_145 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_144 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_143 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_142 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_141 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_140 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_139 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_138 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_137 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_136 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_135 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_134 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_133 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_132 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_131 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_130 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_129 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_128 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_127 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_126 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_125 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_124 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_INHSV6 U1 ( .I(n1), .ZN(n2) );
  LVT_INHSV2SR U2 ( .I(t_m_1_in), .ZN(n1) );
endmodule


module cell_2_3 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
endmodule


module cell_3_123 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_122 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_121 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_120 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_119 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_118 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U5 ( .I(n6), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module cell_3_117 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_116 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_115 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_114 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_113 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_112 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_111 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_110 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_109 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_108 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_107 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_106 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_105 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_104 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_103 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_102 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_101 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_100 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_99 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_98 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_97 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_96 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_95 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8, n9, n10;

  LVT_CLKNHSV0P5 U1 ( .I(t_i_1_in), .ZN(n5) );
  LVT_NAND2HSV2 U2 ( .A1(n8), .A2(n5), .ZN(n6) );
  LVT_NAND2HSV0P5 U3 ( .A1(n4), .A2(t_i_1_in), .ZN(n7) );
  LVT_NAND2HSV2 U4 ( .A1(n6), .A2(n7), .ZN(n9) );
  LVT_INHSV0SR U5 ( .I(n8), .ZN(n4) );
  LVT_NAND2HSV0 U6 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_XOR2HSV2 U7 ( .A1(n10), .A2(n9), .Z(t_i_out) );
  LVT_NAND2HSV0 U8 ( .A1(t_m_1_in), .A2(g_in), .ZN(n10) );
endmodule


module cell_3_94 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_93 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV3 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
  LVT_XNOR2HSV4 U2 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
endmodule


module row_other_3 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1, n2, n3, n4;

  cell_2_3 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_123 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_122 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_121 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_120 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_119 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_118 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_117 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_116 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_115 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_114 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(n4), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_113 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_112 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_111 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_110 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_109 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(n4), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_108 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(n4), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_107 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(n4), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_106 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n4), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_105 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_104 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_103 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_102 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(n2), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_101 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_100 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(n4), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_99 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(n4), 
        .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_98 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_97 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_96 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(n2), 
        .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_95 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_94 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_93 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_CLKNHSV0P5 U1 ( .I(t_m_1_in), .ZN(n3) );
  LVT_INHSV2 U2 ( .I(n3), .ZN(n4) );
  LVT_INHSV0SR U3 ( .I(t_m_1_in), .ZN(n1) );
  LVT_INHSV2 U4 ( .I(n1), .ZN(n2) );
endmodule


module cell_2_2 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_92 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_91 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_90 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_89 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_88 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_87 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_86 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_85 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_84 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_83 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_82 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV2 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_81 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_80 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_79 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_78 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_77 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_76 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_75 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_74 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKXOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_73 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_72 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_71 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_70 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_69 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_68 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_67 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_66 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_65 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_64 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_63 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XNOR2HSV1 U1 ( .A1(n5), .A2(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n2) );
  LVT_NAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_62 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6, n7, n8, n9;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n8) );
  LVT_CLKNAND2HSV2 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n9) );
  LVT_CLKNAND2HSV3 U2 ( .A1(n2), .A2(n4), .ZN(n6) );
  LVT_NAND2HSV0P5 U4 ( .A1(n9), .A2(n7), .ZN(n5) );
  LVT_NAND2HSV4 U5 ( .A1(n5), .A2(n6), .ZN(t_i_out) );
  LVT_INHSV2 U6 ( .I(n9), .ZN(n2) );
  LVT_INHSV2 U7 ( .I(n7), .ZN(n4) );
  LVT_XNOR2HSV4 U8 ( .A1(n8), .A2(t_i_1_in), .ZN(n7) );
endmodule


module row_other_2 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;
  wire   n1;

  cell_2_2 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_92 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_91 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_90 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_89 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_88 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_87 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_86 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_85 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_84 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_83 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_82 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_81 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_80 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_79 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_78 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_77 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_76 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_75 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_74 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_73 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_72 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_71 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_70 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_69 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_68 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_67 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_66 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_65 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_64 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(n1), 
        .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_63 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_62 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
  LVT_BUFHSV2RT U1 ( .I(t_m_1_in), .Z(n1) );
endmodule


module cell_2_1 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4;

  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(n3), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U2 ( .A1(t_m_1_in), .A2(g_in), .ZN(n3) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
endmodule


module cell_3_61 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_60 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_59 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_58 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_57 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_56 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_55 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_54 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_53 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_52 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_51 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_50 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV0P5 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_49 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_48 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_47 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_46 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_45 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_44 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_43 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_42 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_XOR2HSV0 U1 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_CLKNHSV0 U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_41 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_40 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_39 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_38 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_37 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_36 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV4 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
endmodule


module cell_3_35 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_34 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_33 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n5), .A2(n6), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_32 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_31 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n2, n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n5) );
  LVT_CLKNAND2HSV1 U1 ( .A1(n6), .A2(n4), .ZN(n2) );
  LVT_OAI21HSV2 U2 ( .A1(n6), .A2(n4), .B(n2), .ZN(t_i_out) );
  LVT_XNOR2HSV4 U4 ( .A1(t_i_1_in), .A2(n5), .ZN(n4) );
  LVT_CLKNAND2HSV1 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module row_other_1 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_1 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_61 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_60 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_59 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_58 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_57 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_56 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_55 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_54 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_53 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_52 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_51 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_50 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_49 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_48 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_47 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_46 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_45 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_44 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_43 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_42 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_41 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_40 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_39 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_38 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_37 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_36 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_35 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_34 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_33 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_32 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_31 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module cell_2_0 ( a_in, g_in, b_in, t_m_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in;
  output t_i_out;
  wire   n3, n4, n5, n6;

  LVT_OAI21HSV2 U1 ( .A1(n3), .A2(n5), .B(n4), .ZN(t_i_out) );
  LVT_NAND2HSV2 U2 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_NAND2HSV0P5 U3 ( .A1(n3), .A2(n5), .ZN(n4) );
  LVT_CLKNHSV1 U4 ( .I(n6), .ZN(n3) );
  LVT_CLKNAND2HSV1 U5 ( .A1(t_m_1_in), .A2(g_in), .ZN(n5) );
endmodule


module cell_3_30 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV1 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_29 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_28 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_27 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_26 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_NAND2HSV0P5 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_25 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_24 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_23 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_22 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_21 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_20 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_19 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_18 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_17 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_16 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_15 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_14 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_13 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_XOR2HSV0 U2 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_12 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_11 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_10 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_9 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_8 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV1 U1 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U4 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_7 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
endmodule


module cell_3_6 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_5 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_4 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
  LVT_XOR2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
endmodule


module cell_3_3 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_CLKNAND2HSV0 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_XOR2HSV0 U2 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_NAND2HSV2 U5 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U6 ( .I(n6), .ZN(n4) );
endmodule


module cell_3_2 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_1 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6;

  LVT_XOR2HSV0 U2 ( .A1(n4), .A2(t_i_1_in), .Z(n5) );
  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n4) );
  LVT_XOR2HSV0 U1 ( .A1(n6), .A2(n5), .Z(t_i_out) );
  LVT_NAND2HSV0P5 U4 ( .A1(t_m_1_in), .A2(g_in), .ZN(n6) );
endmodule


module cell_3_0 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_out );
  input a_in, g_in, b_in, t_m_1_in, t_i_1_in;
  output t_i_out;
  wire   n4, n5, n6, n7, n8;

  LVT_CLKNAND2HSV0 U3 ( .A1(b_in), .A2(a_in), .ZN(n6) );
  LVT_OAI21HSV2 U1 ( .A1(n4), .A2(t_i_1_in), .B(n5), .ZN(n7) );
  LVT_NAND2HSV2 U2 ( .A1(n4), .A2(t_i_1_in), .ZN(n5) );
  LVT_INHSV0SR U4 ( .I(n6), .ZN(n4) );
  LVT_XOR2HSV0 U5 ( .A1(n8), .A2(n7), .Z(t_i_out) );
  LVT_CLKNAND2HSV1 U6 ( .A1(t_m_1_in), .A2(g_in), .ZN(n8) );
endmodule


module row_other_0 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_out, 
        t_i_2_out );
  input [31:0] a_in;
  input [31:0] g_in;
  input [30:0] t_i_1_in;
  output [30:0] t_i_1_out;
  input b_in, t_m_1_in;
  output t_i_2_out;


  cell_2_0 u0 ( .a_in(a_in[0]), .g_in(g_in[0]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_out(t_i_1_out[0]) );
  cell_3_30 u1 ( .a_in(a_in[1]), .g_in(g_in[1]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[0]), .t_i_out(t_i_1_out[1]) );
  cell_3_29 u2 ( .a_in(a_in[2]), .g_in(g_in[2]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[1]), .t_i_out(t_i_1_out[2]) );
  cell_3_28 u3 ( .a_in(a_in[3]), .g_in(g_in[3]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[2]), .t_i_out(t_i_1_out[3]) );
  cell_3_27 u4 ( .a_in(a_in[4]), .g_in(g_in[4]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[3]), .t_i_out(t_i_1_out[4]) );
  cell_3_26 u5 ( .a_in(a_in[5]), .g_in(g_in[5]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[4]), .t_i_out(t_i_1_out[5]) );
  cell_3_25 u6 ( .a_in(a_in[6]), .g_in(g_in[6]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[5]), .t_i_out(t_i_1_out[6]) );
  cell_3_24 u7 ( .a_in(a_in[7]), .g_in(g_in[7]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[6]), .t_i_out(t_i_1_out[7]) );
  cell_3_23 u8 ( .a_in(a_in[8]), .g_in(g_in[8]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[7]), .t_i_out(t_i_1_out[8]) );
  cell_3_22 u9 ( .a_in(a_in[9]), .g_in(g_in[9]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[8]), .t_i_out(t_i_1_out[9]) );
  cell_3_21 u10 ( .a_in(a_in[10]), .g_in(g_in[10]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[9]), .t_i_out(t_i_1_out[10]) );
  cell_3_20 u11 ( .a_in(a_in[11]), .g_in(g_in[11]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[10]), .t_i_out(t_i_1_out[11]) );
  cell_3_19 u12 ( .a_in(a_in[12]), .g_in(g_in[12]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[11]), .t_i_out(t_i_1_out[12]) );
  cell_3_18 u13 ( .a_in(a_in[13]), .g_in(g_in[13]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[12]), .t_i_out(t_i_1_out[13]) );
  cell_3_17 u14 ( .a_in(a_in[14]), .g_in(g_in[14]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[13]), .t_i_out(t_i_1_out[14]) );
  cell_3_16 u15 ( .a_in(a_in[15]), .g_in(g_in[15]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[14]), .t_i_out(t_i_1_out[15]) );
  cell_3_15 u16 ( .a_in(a_in[16]), .g_in(g_in[16]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[15]), .t_i_out(t_i_1_out[16]) );
  cell_3_14 u17 ( .a_in(a_in[17]), .g_in(g_in[17]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[16]), .t_i_out(t_i_1_out[17]) );
  cell_3_13 u18 ( .a_in(a_in[18]), .g_in(g_in[18]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[17]), .t_i_out(t_i_1_out[18]) );
  cell_3_12 u19 ( .a_in(a_in[19]), .g_in(g_in[19]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[18]), .t_i_out(t_i_1_out[19]) );
  cell_3_11 u20 ( .a_in(a_in[20]), .g_in(g_in[20]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[19]), .t_i_out(t_i_1_out[20]) );
  cell_3_10 u21 ( .a_in(a_in[21]), .g_in(g_in[21]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[20]), .t_i_out(t_i_1_out[21]) );
  cell_3_9 u22 ( .a_in(a_in[22]), .g_in(g_in[22]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[21]), .t_i_out(t_i_1_out[22]) );
  cell_3_8 u23 ( .a_in(a_in[23]), .g_in(g_in[23]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[22]), .t_i_out(t_i_1_out[23]) );
  cell_3_7 u24 ( .a_in(a_in[24]), .g_in(g_in[24]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[23]), .t_i_out(t_i_1_out[24]) );
  cell_3_6 u25 ( .a_in(a_in[25]), .g_in(g_in[25]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[24]), .t_i_out(t_i_1_out[25]) );
  cell_3_5 u26 ( .a_in(a_in[26]), .g_in(g_in[26]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[25]), .t_i_out(t_i_1_out[26]) );
  cell_3_4 u27 ( .a_in(a_in[27]), .g_in(g_in[27]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[26]), .t_i_out(t_i_1_out[27]) );
  cell_3_3 u28 ( .a_in(a_in[28]), .g_in(g_in[28]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[27]), .t_i_out(t_i_1_out[28]) );
  cell_3_2 u29 ( .a_in(a_in[29]), .g_in(g_in[29]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[28]), .t_i_out(t_i_1_out[29]) );
  cell_3_1 u30 ( .a_in(a_in[30]), .g_in(g_in[30]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[29]), .t_i_out(t_i_1_out[30]) );
  cell_3_0 u31 ( .a_in(a_in[31]), .g_in(g_in[31]), .b_in(b_in), .t_m_1_in(
        t_m_1_in), .t_i_1_in(t_i_1_in[30]), .t_i_out(t_i_2_out) );
endmodule


module PE_core_0 ( a_in, g_in, b_in, t_m_1_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, t_i_1_out, t_i_2_out, t_i_1_out_0 );
  input [31:0] a_in;
  input [31:0] g_in;
  input [31:0] b_in;
  input [31:0] t_m_1_in;
  input [30:0] t_i_1_in;
  input [30:0] t_i_2_in;
  output [31:0] a_out;
  output [31:0] g_out;
  output [30:0] t_i_1_out;
  output [30:0] t_i_2_out;
  input t_i_1_in_0;
  output t_i_1_out_0;
  wire   n1, n2, n4, n6, n7, n9, n10, n12, n13, n15, n16, n18, n21, n23, n24;
  wire   [30:0] t0;
  wire   [30:0] t1;
  wire   [30:0] t2;
  wire   [30:0] t3;
  wire   [30:0] t4;
  wire   [30:0] t5;
  wire   [30:0] t6;
  wire   [30:0] t7;
  wire   [30:0] t8;
  wire   [30:0] t9;
  wire   [30:0] t10;
  wire   [30:0] t11;
  wire   [30:0] t12;
  wire   [30:0] t13;
  wire   [30:0] t14;
  wire   [30:0] t15;
  wire   [30:0] t16;
  wire   [30:0] t17;
  wire   [30:0] t18;
  wire   [30:0] t19;
  wire   [30:0] t20;
  wire   [30:0] t21;
  wire   [30:0] t22;
  wire   [30:0] t23;
  wire   [30:0] t24;
  wire   [30:0] t25;
  wire   [30:0] t26;
  wire   [30:0] t27;
  wire   [30:0] t28;
  wire   [30:0] t29;
  wire   [30:0] t30;
  assign a_out[29] = a_in[29];
  assign a_out[27] = a_in[27];
  assign a_out[26] = a_in[26];
  assign a_out[22] = a_in[22];
  assign a_out[20] = a_in[20];
  assign a_out[19] = a_in[19];
  assign a_out[18] = a_in[18];
  assign a_out[17] = a_in[17];
  assign a_out[16] = a_in[16];
  assign a_out[15] = a_in[15];
  assign a_out[14] = a_in[14];
  assign a_out[13] = a_in[13];
  assign a_out[12] = a_in[12];
  assign a_out[11] = a_in[11];
  assign a_out[10] = a_in[10];
  assign a_out[9] = a_in[9];
  assign a_out[8] = a_in[8];
  assign a_out[7] = a_in[7];
  assign a_out[6] = a_in[6];
  assign a_out[5] = a_in[5];
  assign a_out[4] = a_in[4];
  assign a_out[3] = a_in[3];
  assign a_out[2] = a_in[2];
  assign a_out[1] = a_in[1];
  assign a_out[0] = a_in[0];
  assign g_out[31] = g_in[31];
  assign g_out[30] = g_in[30];
  assign g_out[29] = g_in[29];
  assign g_out[28] = g_in[28];
  assign g_out[27] = g_in[27];
  assign g_out[25] = g_in[25];
  assign g_out[24] = g_in[24];
  assign g_out[22] = g_in[22];
  assign g_out[21] = g_in[21];
  assign g_out[20] = g_in[20];
  assign g_out[19] = g_in[19];
  assign g_out[18] = g_in[18];
  assign g_out[17] = g_in[17];
  assign g_out[16] = g_in[16];
  assign g_out[15] = g_in[15];
  assign g_out[14] = g_in[14];
  assign g_out[13] = g_in[13];
  assign g_out[12] = g_in[12];
  assign g_out[11] = g_in[11];
  assign g_out[10] = g_in[10];
  assign g_out[9] = g_in[9];
  assign g_out[8] = g_in[8];
  assign g_out[7] = g_in[7];
  assign g_out[6] = g_in[6];
  assign g_out[5] = g_in[5];
  assign g_out[4] = g_in[4];
  assign g_out[3] = g_in[3];
  assign g_out[2] = g_in[2];
  assign g_out[1] = g_in[1];
  assign g_out[0] = g_in[0];

  row_1_0 u0 ( .a_in({n24, a_in[30:29], n13, a_in[27:25], n16, n7, a_in[22], 
        n4, a_in[20:0]}), .g_in({g_in[31:27], n2, g_in[25:24], n10, g_in[22:0]}), .b_in(b_in[31]), .t_m_1_in(t_m_1_in[31]), .t_i_1_in({t_i_1_in, t_i_1_in_0}), 
        .t_i_2_in(t_i_2_in), .t_i_1_out(t0), .t_i_2_out(t_i_2_out[30]) );
  row_other_30 u1 ( .a_in({n24, a_out[30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[30]), 
        .t_m_1_in(t_m_1_in[30]), .t_i_1_in(t0), .t_i_1_out(t1), .t_i_2_out(
        t_i_2_out[29]) );
  row_other_29 u2 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[29]), 
        .t_m_1_in(t_m_1_in[29]), .t_i_1_in(t1), .t_i_1_out(t2), .t_i_2_out(
        t_i_2_out[28]) );
  row_other_28 u3 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[28]), 
        .t_m_1_in(t_m_1_in[28]), .t_i_1_in(t2), .t_i_1_out(t3), .t_i_2_out(
        t_i_2_out[27]) );
  row_other_27 u4 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[27]), 
        .t_m_1_in(t_m_1_in[27]), .t_i_1_in(t3), .t_i_1_out(t4), .t_i_2_out(
        t_i_2_out[26]) );
  row_other_26 u5 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[26]), 
        .t_m_1_in(t_m_1_in[26]), .t_i_1_in(t4), .t_i_1_out(t5), .t_i_2_out(
        t_i_2_out[25]) );
  row_other_25 u6 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[25]), 
        .t_m_1_in(t_m_1_in[25]), .t_i_1_in(t5), .t_i_1_out(t6), .t_i_2_out(
        t_i_2_out[24]) );
  row_other_24 u7 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[24]), 
        .t_m_1_in(t_m_1_in[24]), .t_i_1_in(t6), .t_i_1_out(t7), .t_i_2_out(
        t_i_2_out[23]) );
  row_other_23 u8 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[23]), 
        .t_m_1_in(t_m_1_in[23]), .t_i_1_in(t7), .t_i_1_out(t8), .t_i_2_out(
        t_i_2_out[22]) );
  row_other_22 u9 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[22]), 
        .t_m_1_in(t_m_1_in[22]), .t_i_1_in(t8), .t_i_1_out(t9), .t_i_2_out(
        t_i_2_out[21]) );
  row_other_21 u10 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[21]), 
        .t_m_1_in(t_m_1_in[21]), .t_i_1_in(t9), .t_i_1_out(t10), .t_i_2_out(
        t_i_2_out[20]) );
  row_other_20 u11 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[20]), 
        .t_m_1_in(t_m_1_in[20]), .t_i_1_in(t10), .t_i_1_out(t11), .t_i_2_out(
        t_i_2_out[19]) );
  row_other_19 u12 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[19]), 
        .t_m_1_in(t_m_1_in[19]), .t_i_1_in(t11), .t_i_1_out(t12), .t_i_2_out(
        t_i_2_out[18]) );
  row_other_18 u13 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[18]), 
        .t_m_1_in(t_m_1_in[18]), .t_i_1_in(t12), .t_i_1_out(t13), .t_i_2_out(
        t_i_2_out[17]) );
  row_other_17 u14 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[17]), 
        .t_m_1_in(t_m_1_in[17]), .t_i_1_in(t13), .t_i_1_out(t14), .t_i_2_out(
        t_i_2_out[16]) );
  row_other_16 u15 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[16]), 
        .t_m_1_in(t_m_1_in[16]), .t_i_1_in(t14), .t_i_1_out(t15), .t_i_2_out(
        t_i_2_out[15]) );
  row_other_15 u16 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[15]), 
        .t_m_1_in(t_m_1_in[15]), .t_i_1_in(t15), .t_i_1_out(t16), .t_i_2_out(
        t_i_2_out[14]) );
  row_other_14 u17 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[14]), 
        .t_m_1_in(t_m_1_in[14]), .t_i_1_in(t16), .t_i_1_out(t17), .t_i_2_out(
        t_i_2_out[13]) );
  row_other_13 u18 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[13]), 
        .t_m_1_in(t_m_1_in[13]), .t_i_1_in(t17), .t_i_1_out(t18), .t_i_2_out(
        t_i_2_out[12]) );
  row_other_12 u19 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[12]), 
        .t_m_1_in(t_m_1_in[12]), .t_i_1_in(t18), .t_i_1_out(t19), .t_i_2_out(
        t_i_2_out[11]) );
  row_other_11 u20 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[11]), 
        .t_m_1_in(t_m_1_in[11]), .t_i_1_in(t19), .t_i_1_out(t20), .t_i_2_out(
        t_i_2_out[10]) );
  row_other_10 u21 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[10]), 
        .t_m_1_in(t_m_1_in[10]), .t_i_1_in(t20), .t_i_1_out(t21), .t_i_2_out(
        t_i_2_out[9]) );
  row_other_9 u22 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[9]), 
        .t_m_1_in(t_m_1_in[9]), .t_i_1_in(t21), .t_i_1_out(t22), .t_i_2_out(
        t_i_2_out[8]) );
  row_other_8 u23 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[8]), 
        .t_m_1_in(t_m_1_in[8]), .t_i_1_in(t22), .t_i_1_out(t23), .t_i_2_out(
        t_i_2_out[7]) );
  row_other_7 u24 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[7]), 
        .t_m_1_in(t_m_1_in[7]), .t_i_1_in(t23), .t_i_1_out(t24), .t_i_2_out(
        t_i_2_out[6]) );
  row_other_6 u25 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[6]), 
        .t_m_1_in(t_m_1_in[6]), .t_i_1_in(t24), .t_i_1_out(t25), .t_i_2_out(
        t_i_2_out[5]) );
  row_other_5 u26 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[5]), 
        .t_m_1_in(t_m_1_in[5]), .t_i_1_in(t25), .t_i_1_out(t26), .t_i_2_out(
        t_i_2_out[4]) );
  row_other_4 u27 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[4]), 
        .t_m_1_in(t_m_1_in[4]), .t_i_1_in(t26), .t_i_1_out(t27), .t_i_2_out(
        t_i_2_out[3]) );
  row_other_3 u28 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[3]), 
        .t_m_1_in(t_m_1_in[3]), .t_i_1_in(t27), .t_i_1_out(t28), .t_i_2_out(
        t_i_2_out[2]) );
  row_other_2 u29 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[2]), 
        .t_m_1_in(t_m_1_in[2]), .t_i_1_in(t28), .t_i_1_out(t29), .t_i_2_out(
        t_i_2_out[1]) );
  row_other_1 u30 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[1]), 
        .t_m_1_in(t_m_1_in[1]), .t_i_1_in(t29), .t_i_1_out(t30), .t_i_2_out(
        t_i_2_out[0]) );
  row_other_0 u31 ( .a_in({a_out[31:30], a_in[29], a_out[28], a_in[27:26], 
        a_out[25:23], a_in[22], a_out[21], a_in[20:0]}), .g_in({g_in[31:27], 
        g_out[26], g_in[25:24], g_out[23], g_in[22:0]}), .b_in(b_in[0]), 
        .t_m_1_in(t_m_1_in[0]), .t_i_1_in(t30), .t_i_1_out(t_i_1_out), 
        .t_i_2_out(t_i_1_out_0) );
  LVT_INHSV3SR U1 ( .I(g_in[26]), .ZN(n1) );
  LVT_CLKNHSV2P5 U2 ( .I(n1), .ZN(n2) );
  LVT_INHSV2SR U3 ( .I(n1), .ZN(g_out[26]) );
  LVT_INHSV2 U4 ( .I(n9), .ZN(n10) );
  LVT_INHSV2 U5 ( .I(a_in[23]), .ZN(n6) );
  LVT_INHSV2 U6 ( .I(a_in[24]), .ZN(n15) );
  LVT_INHSV2 U7 ( .I(a_in[28]), .ZN(n12) );
  LVT_INHSV2 U8 ( .I(g_in[23]), .ZN(n9) );
  LVT_BUFHSV2 U9 ( .I(a_in[21]), .Z(n4) );
  LVT_BUFHSV2RT U10 ( .I(a_in[21]), .Z(a_out[21]) );
  LVT_INHSV2SR U11 ( .I(n6), .ZN(n7) );
  LVT_INHSV2SR U12 ( .I(n6), .ZN(a_out[23]) );
  LVT_INHSV2SR U13 ( .I(n9), .ZN(g_out[23]) );
  LVT_INHSV2SR U14 ( .I(n12), .ZN(n13) );
  LVT_INHSV2SR U15 ( .I(n12), .ZN(a_out[28]) );
  LVT_CLKNHSV2 U16 ( .I(n15), .ZN(n16) );
  LVT_INHSV2SR U17 ( .I(n15), .ZN(a_out[24]) );
  LVT_INHSV2 U18 ( .I(a_in[25]), .ZN(n18) );
  LVT_INHSV2SR U19 ( .I(n18), .ZN(a_out[25]) );
  LVT_INHSV2 U20 ( .I(a_in[31]), .ZN(n23) );
  LVT_INHSV2 U21 ( .I(n23), .ZN(n24) );
  LVT_INHSV2 U22 ( .I(a_in[30]), .ZN(n21) );
  LVT_BUFHSV2 U23 ( .I(a_in[31]), .Z(a_out[31]) );
  LVT_CLKNHSV2 U24 ( .I(n21), .ZN(a_out[30]) );
endmodule


module regist_32bit_1 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n2), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n2), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n2), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_32bit_0 ( clk, rstn, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV1 \out_reg[31]  ( .D(in[31]), .CK(clk), .RDN(n1), .Q(out[31]) );
  LVT_DRNQHSV1 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV1 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV1 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV1 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV1 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV1 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV1 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV1 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV1 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV1 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV1 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV1 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV1 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV1 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV1 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV1 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV1 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV1 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV1 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV1 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV1 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV1 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV1 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV1 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(n2), .Q(out[7]) );
  LVT_DRNQHSV1 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n1), .Q(out[6]) );
  LVT_DRNQHSV1 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n2), .Q(out[5]) );
  LVT_DRNQHSV1 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n1), .Q(out[4]) );
  LVT_DRNQHSV1 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n2), .Q(out[3]) );
  LVT_DRNQHSV1 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n1), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n2), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module regist_31bit_0 ( clk, rstn, in, out );
  input [30:0] in;
  output [30:0] out;
  input clk, rstn;
  wire   n1, n2, n3;

  LVT_DRNQHSV2 \out_reg[30]  ( .D(in[30]), .CK(clk), .RDN(n1), .Q(out[30]) );
  LVT_DRNQHSV2 \out_reg[29]  ( .D(in[29]), .CK(clk), .RDN(n1), .Q(out[29]) );
  LVT_DRNQHSV2 \out_reg[28]  ( .D(in[28]), .CK(clk), .RDN(n1), .Q(out[28]) );
  LVT_DRNQHSV2 \out_reg[27]  ( .D(in[27]), .CK(clk), .RDN(n1), .Q(out[27]) );
  LVT_DRNQHSV2 \out_reg[26]  ( .D(in[26]), .CK(clk), .RDN(n1), .Q(out[26]) );
  LVT_DRNQHSV2 \out_reg[25]  ( .D(in[25]), .CK(clk), .RDN(n1), .Q(out[25]) );
  LVT_DRNQHSV2 \out_reg[24]  ( .D(in[24]), .CK(clk), .RDN(n1), .Q(out[24]) );
  LVT_DRNQHSV2 \out_reg[23]  ( .D(in[23]), .CK(clk), .RDN(n1), .Q(out[23]) );
  LVT_DRNQHSV2 \out_reg[22]  ( .D(in[22]), .CK(clk), .RDN(n1), .Q(out[22]) );
  LVT_DRNQHSV2 \out_reg[21]  ( .D(in[21]), .CK(clk), .RDN(n1), .Q(out[21]) );
  LVT_DRNQHSV2 \out_reg[20]  ( .D(in[20]), .CK(clk), .RDN(n1), .Q(out[20]) );
  LVT_DRNQHSV2 \out_reg[19]  ( .D(in[19]), .CK(clk), .RDN(n2), .Q(out[19]) );
  LVT_DRNQHSV2 \out_reg[18]  ( .D(in[18]), .CK(clk), .RDN(n2), .Q(out[18]) );
  LVT_DRNQHSV2 \out_reg[17]  ( .D(in[17]), .CK(clk), .RDN(n2), .Q(out[17]) );
  LVT_DRNQHSV2 \out_reg[16]  ( .D(in[16]), .CK(clk), .RDN(n2), .Q(out[16]) );
  LVT_DRNQHSV2 \out_reg[15]  ( .D(in[15]), .CK(clk), .RDN(n2), .Q(out[15]) );
  LVT_DRNQHSV2 \out_reg[14]  ( .D(in[14]), .CK(clk), .RDN(n2), .Q(out[14]) );
  LVT_DRNQHSV2 \out_reg[13]  ( .D(in[13]), .CK(clk), .RDN(n2), .Q(out[13]) );
  LVT_DRNQHSV2 \out_reg[12]  ( .D(in[12]), .CK(clk), .RDN(n2), .Q(out[12]) );
  LVT_DRNQHSV2 \out_reg[11]  ( .D(in[11]), .CK(clk), .RDN(n2), .Q(out[11]) );
  LVT_DRNQHSV2 \out_reg[10]  ( .D(in[10]), .CK(clk), .RDN(n2), .Q(out[10]) );
  LVT_DRNQHSV2 \out_reg[9]  ( .D(in[9]), .CK(clk), .RDN(n2), .Q(out[9]) );
  LVT_DRNQHSV2 \out_reg[8]  ( .D(in[8]), .CK(clk), .RDN(n2), .Q(out[8]) );
  LVT_DRNQHSV2 \out_reg[7]  ( .D(in[7]), .CK(clk), .RDN(rstn), .Q(out[7]) );
  LVT_DRNQHSV2 \out_reg[6]  ( .D(in[6]), .CK(clk), .RDN(n2), .Q(out[6]) );
  LVT_DRNQHSV2 \out_reg[5]  ( .D(in[5]), .CK(clk), .RDN(n1), .Q(out[5]) );
  LVT_DRNQHSV2 \out_reg[4]  ( .D(in[4]), .CK(clk), .RDN(n2), .Q(out[4]) );
  LVT_DRNQHSV2 \out_reg[3]  ( .D(in[3]), .CK(clk), .RDN(n1), .Q(out[3]) );
  LVT_DRNQHSV2 \out_reg[2]  ( .D(in[2]), .CK(clk), .RDN(n2), .Q(out[2]) );
  LVT_DRNQHSV2 \out_reg[1]  ( .D(in[1]), .CK(clk), .RDN(n1), .Q(out[1]) );
  LVT_DRNQHSV2 \out_reg[0]  ( .D(in[0]), .CK(clk), .RDN(n1), .Q(out[0]) );
  LVT_INHSV2 U3 ( .I(rstn), .ZN(n3) );
  LVT_INHSV2 U4 ( .I(n3), .ZN(n2) );
  LVT_INHSV2 U5 ( .I(n3), .ZN(n1) );
endmodule


module PE_0 ( clk, rstn, ctr, a_in, g_in, b_in, t_i_1_in, t_i_1_in_0, t_i_2_in, 
        a_out, g_out, b_out, t_i_1_out, t_i_2_out, t_i_1_out_0, ctro );
  input [31:0] a_in;
  input [31:0] g_in;
  input [31:0] b_in;
  input [30:0] t_i_1_in;
  input [30:0] t_i_2_in;
  output [31:0] a_out;
  output [31:0] g_out;
  output [31:0] b_out;
  output [30:0] t_i_1_out;
  output [30:0] t_i_2_out;
  input clk, rstn, ctr, t_i_1_in_0;
  output t_i_1_out_0, ctro;
  wire   n109, n110, n111, l_ctr, l_t_i_1_in_0, \c_t_i_1_in[0] , c_t_i_1_in_0,
         to_1, ti_1, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n35, n36, n37, n38, n39,
         n40, n41, n42, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108;
  wire   [31:0] l_a;
  wire   [31:0] l_g;
  wire   [30:0] l_t_i_1_in;
  wire   [30:0] l_t_i_2_in;
  wire   [31:0] mux_b;
  wire   [31:0] mux_bq;
  wire   [30:0] to_7;
  wire   [30:0] ti_7;
  wire   [31:0] ao;
  wire   [31:0] go;
  wire   [30:0] to;

  LVT_AO22HSV0 U35 ( .A1(mux_bq[9]), .A2(n41), .B1(b_out[9]), .B2(n106), .Z(
        mux_b[9]) );
  LVT_AO22HSV0 U36 ( .A1(mux_bq[8]), .A2(n41), .B1(b_out[8]), .B2(n106), .Z(
        mux_b[8]) );
  LVT_AO22HSV0 U37 ( .A1(mux_bq[7]), .A2(n41), .B1(b_out[7]), .B2(n106), .Z(
        mux_b[7]) );
  LVT_AO22HSV0 U38 ( .A1(mux_bq[6]), .A2(n41), .B1(b_out[6]), .B2(n106), .Z(
        mux_b[6]) );
  LVT_AO22HSV0 U39 ( .A1(mux_bq[5]), .A2(n41), .B1(b_out[5]), .B2(n106), .Z(
        mux_b[5]) );
  LVT_AO22HSV0 U40 ( .A1(mux_bq[4]), .A2(n41), .B1(b_out[4]), .B2(n106), .Z(
        mux_b[4]) );
  LVT_AO22HSV0 U41 ( .A1(mux_bq[3]), .A2(n41), .B1(b_out[3]), .B2(n106), .Z(
        mux_b[3]) );
  LVT_AO22HSV0 U42 ( .A1(n21), .A2(n41), .B1(b_out[31]), .B2(n106), .Z(
        mux_b[31]) );
  LVT_AO22HSV0 U43 ( .A1(mux_bq[30]), .A2(n41), .B1(b_out[30]), .B2(n106), .Z(
        mux_b[30]) );
  LVT_AO22HSV0 U44 ( .A1(mux_bq[2]), .A2(n41), .B1(b_out[2]), .B2(n106), .Z(
        mux_b[2]) );
  LVT_AO22HSV0 U45 ( .A1(mux_bq[29]), .A2(n41), .B1(b_out[29]), .B2(n106), .Z(
        mux_b[29]) );
  LVT_AO22HSV0 U46 ( .A1(mux_bq[28]), .A2(n41), .B1(b_out[28]), .B2(n106), .Z(
        mux_b[28]) );
  LVT_AO22HSV0 U47 ( .A1(mux_bq[27]), .A2(n41), .B1(b_out[27]), .B2(n106), .Z(
        mux_b[27]) );
  LVT_AO22HSV0 U48 ( .A1(mux_bq[26]), .A2(n41), .B1(b_out[26]), .B2(n106), .Z(
        mux_b[26]) );
  LVT_AO22HSV0 U49 ( .A1(mux_bq[25]), .A2(n41), .B1(b_out[25]), .B2(n106), .Z(
        mux_b[25]) );
  LVT_AO22HSV0 U50 ( .A1(mux_bq[24]), .A2(n41), .B1(b_out[24]), .B2(n106), .Z(
        mux_b[24]) );
  LVT_AO22HSV0 U51 ( .A1(mux_bq[23]), .A2(n41), .B1(b_out[23]), .B2(n106), .Z(
        mux_b[23]) );
  LVT_AO22HSV0 U52 ( .A1(mux_bq[22]), .A2(n41), .B1(b_out[22]), .B2(n106), .Z(
        mux_b[22]) );
  LVT_AO22HSV0 U53 ( .A1(mux_bq[21]), .A2(n41), .B1(b_out[21]), .B2(n106), .Z(
        mux_b[21]) );
  LVT_AO22HSV0 U54 ( .A1(mux_bq[20]), .A2(n41), .B1(b_out[20]), .B2(n106), .Z(
        mux_b[20]) );
  LVT_AO22HSV0 U55 ( .A1(mux_bq[1]), .A2(n41), .B1(b_out[1]), .B2(n106), .Z(
        mux_b[1]) );
  LVT_AO22HSV0 U56 ( .A1(mux_bq[19]), .A2(n41), .B1(b_out[19]), .B2(n106), .Z(
        mux_b[19]) );
  LVT_AO22HSV0 U57 ( .A1(mux_bq[18]), .A2(n41), .B1(b_out[18]), .B2(n106), .Z(
        mux_b[18]) );
  LVT_AO22HSV0 U58 ( .A1(mux_bq[17]), .A2(n41), .B1(b_out[17]), .B2(n106), .Z(
        mux_b[17]) );
  LVT_AO22HSV0 U59 ( .A1(mux_bq[16]), .A2(n41), .B1(b_out[16]), .B2(n106), .Z(
        mux_b[16]) );
  LVT_AO22HSV0 U60 ( .A1(mux_bq[15]), .A2(n41), .B1(b_out[15]), .B2(n106), .Z(
        mux_b[15]) );
  LVT_AO22HSV0 U61 ( .A1(mux_bq[14]), .A2(n41), .B1(b_out[14]), .B2(n106), .Z(
        mux_b[14]) );
  LVT_AO22HSV0 U62 ( .A1(mux_bq[13]), .A2(n41), .B1(b_out[13]), .B2(n106), .Z(
        mux_b[13]) );
  LVT_AO22HSV0 U63 ( .A1(mux_bq[12]), .A2(n41), .B1(b_out[12]), .B2(n106), .Z(
        mux_b[12]) );
  LVT_AO22HSV0 U64 ( .A1(mux_bq[11]), .A2(n41), .B1(b_out[11]), .B2(n106), .Z(
        mux_b[11]) );
  LVT_AO22HSV0 U65 ( .A1(mux_bq[10]), .A2(n41), .B1(b_out[10]), .B2(n106), .Z(
        mux_b[10]) );
  LVT_AO22HSV0 U66 ( .A1(mux_bq[0]), .A2(n41), .B1(b_out[0]), .B2(n106), .Z(
        mux_b[0]) );
  LVT_NOR2HSV0 U67 ( .A1(n107), .A2(n106), .ZN(c_t_i_1_in_0) );
  LVT_AOI21HSV0 U69 ( .A1(n105), .A2(n104), .B(n106), .ZN(\c_t_i_1_in[0] ) );
  LVT_AND4HSV0 U71 ( .A1(n103), .A2(n102), .A3(n101), .A4(n100), .Z(n104) );
  LVT_NOR4HSV0 U72 ( .A1(l_t_i_1_in[9]), .A2(l_t_i_1_in[8]), .A3(l_t_i_1_in[7]), .A4(l_t_i_1_in[6]), .ZN(n100) );
  LVT_NOR4HSV0 U73 ( .A1(l_t_i_1_in[5]), .A2(l_t_i_1_in[4]), .A3(l_t_i_1_in[3]), .A4(l_t_i_1_in[30]), .ZN(n101) );
  LVT_NOR4HSV0 U74 ( .A1(l_t_i_1_in[2]), .A2(l_t_i_1_in[29]), .A3(
        l_t_i_1_in[28]), .A4(l_t_i_1_in[27]), .ZN(n102) );
  LVT_NOR4HSV0 U75 ( .A1(l_t_i_1_in[26]), .A2(l_t_i_1_in[25]), .A3(
        l_t_i_1_in[24]), .A4(l_t_i_1_in[23]), .ZN(n103) );
  LVT_AND4HSV0 U76 ( .A1(n99), .A2(n98), .A3(n97), .A4(n96), .Z(n105) );
  LVT_NOR4HSV0 U77 ( .A1(l_t_i_1_in[22]), .A2(l_t_i_1_in[21]), .A3(
        l_t_i_1_in[20]), .A4(l_t_i_1_in[1]), .ZN(n96) );
  LVT_NOR4HSV0 U78 ( .A1(l_t_i_1_in[19]), .A2(l_t_i_1_in[18]), .A3(
        l_t_i_1_in[17]), .A4(l_t_i_1_in[16]), .ZN(n97) );
  LVT_NOR4HSV0 U79 ( .A1(l_t_i_1_in[15]), .A2(l_t_i_1_in[14]), .A3(
        l_t_i_1_in[13]), .A4(l_t_i_1_in[12]), .ZN(n98) );
  LVT_NOR3HSV0 U80 ( .A1(l_t_i_1_in[0]), .A2(l_t_i_1_in[11]), .A3(
        l_t_i_1_in[10]), .ZN(n99) );
  regist_32bit_5 u0 ( .clk(clk), .rstn(n94), .in(a_in), .out(l_a) );
  regist_32bit_4 u1 ( .clk(clk), .rstn(n94), .in(b_in), .out(b_out) );
  regist_32bit_3 u2 ( .clk(clk), .rstn(n94), .in(g_in), .out(l_g) );
  regist_1bit_3 u3 ( .clk(clk), .rstn(n94), .in(ctr), .out(l_ctr) );
  regist_1bit_2 u4 ( .clk(clk), .rstn(n94), .in(n41), .out(n111) );
  regist_31bit_3 u5 ( .clk(clk), .rstn(n94), .in(t_i_1_in), .out(l_t_i_1_in)
         );
  regist_31bit_2 u6 ( .clk(clk), .rstn(n94), .in(t_i_2_in), .out(l_t_i_2_in)
         );
  regist_1bit_1 u7 ( .clk(clk), .rstn(n94), .in(t_i_1_in_0), .out(l_t_i_1_in_0) );
  regist_32bit_2 u9 ( .clk(clk), .rstn(n94), .in(mux_b), .out(mux_bq) );
  regist_1bit_0 u10 ( .clk(clk), .rstn(n94), .in(to_1), .out(ti_1) );
  regist_31bit_1 u11 ( .clk(clk), .rstn(n94), .in({to_7[30], n72, n73, n67, 
        n66, to_7[25:21], n27, to_7[19], n78, n79, n25, to_7[15:14], n80, n81, 
        n23, n82, n74, n75, to_7[7], n29, to_7[5], n32, to_7[3], n76, to_7[1], 
        n77}), .out(ti_7) );
  PE_core_0 pe ( .a_in(l_a), .g_in({n31, l_g[30:0]}), .b_in({n21, mux_bq[30:0]}), .t_m_1_in({to_1, to_7[30], n72, n73, n67, n66, to_7[25:21], n27, to_7[19], 
        n78, n79, n25, to_7[15:14], n80, n81, n23, n82, n74, n75, to_7[7], n29, 
        to_7[5], n32, to_7[3], n76, to_7[1], n77}), .t_i_1_in({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, \c_t_i_1_in[0] }), .t_i_1_in_0(c_t_i_1_in_0), 
        .t_i_2_in(l_t_i_2_in), .a_out(ao), .g_out(go), .t_i_1_out(to), 
        .t_i_2_out({t_i_2_out[30:17], n109, t_i_2_out[15:3], n110, 
        t_i_2_out[1:0]}), .t_i_1_out_0(t_i_1_out_0) );
  regist_32bit_1 u12 ( .clk(clk), .rstn(n94), .in(ao), .out(a_out) );
  regist_32bit_0 u13 ( .clk(clk), .rstn(n94), .in(go), .out(g_out) );
  regist_31bit_0 u14 ( .clk(clk), .rstn(n94), .in(to), .out(t_i_1_out) );
  LVT_INHSV10 U2 ( .I(n57), .ZN(n77) );
  LVT_INHSV6 U3 ( .I(n64), .ZN(n82) );
  LVT_CLKNHSV5 U4 ( .I(n68), .ZN(n78) );
  LVT_INHSV10 U5 ( .I(n24), .ZN(n25) );
  LVT_CLKNAND2HSV3 U6 ( .A1(t_i_2_out[6]), .A2(n108), .ZN(n17) );
  LVT_CLKNAND2HSV2 U7 ( .A1(t_i_2_out[23]), .A2(n108), .ZN(n37) );
  LVT_IAO22HSV4 U8 ( .B1(t_i_2_out[27]), .B2(n108), .A1(n46), .A2(n108), .ZN(
        n45) );
  LVT_INHSV6 U9 ( .I(n40), .ZN(n66) );
  LVT_INHSV4SR U10 ( .I(n65), .ZN(n75) );
  LVT_AND2HSV4 U11 ( .A1(t_i_2_out[14]), .A2(n108), .Z(n90) );
  LVT_INHSV6SR U12 ( .I(n70), .ZN(n80) );
  LVT_CLKNAND2HSV3 U13 ( .A1(t_i_2_out[30]), .A2(n108), .ZN(n86) );
  LVT_INHSV12 U14 ( .I(n28), .ZN(n29) );
  LVT_NAND2HSV8 U15 ( .A1(n86), .A2(n85), .ZN(to_7[30]) );
  LVT_CLKNHSV8 U16 ( .I(l_ctr), .ZN(n93) );
  LVT_CLKNAND2HSV4 U17 ( .A1(n56), .A2(n55), .ZN(to_7[7]) );
  LVT_NAND2HSV4 U18 ( .A1(t_i_2_out[7]), .A2(n108), .ZN(n56) );
  LVT_INHSV2 U19 ( .I(n44), .ZN(n81) );
  LVT_CLKNAND2HSV4 U20 ( .A1(n37), .A2(n33), .ZN(to_7[23]) );
  LVT_OR2HSV16RD U21 ( .A1(n90), .A2(n89), .Z(to_7[14]) );
  LVT_NAND2HSV3 U22 ( .A1(ti_1), .A2(l_ctr), .ZN(n91) );
  LVT_AOI22HSV2 U23 ( .A1(ti_7[12]), .A2(n111), .B1(t_i_2_out[12]), .B2(n108), 
        .ZN(n44) );
  LVT_INHSV10SR U24 ( .I(n71), .ZN(n72) );
  LVT_CLKNAND2HSV8 U25 ( .A1(l_t_i_1_in_0), .A2(n93), .ZN(n92) );
  LVT_INHSV12SR U26 ( .I(n26), .ZN(n27) );
  LVT_CLKNAND2HSV8 U27 ( .A1(n53), .A2(n54), .ZN(to_7[24]) );
  LVT_NAND2HSV0P5 U28 ( .A1(t_i_2_out[11]), .A2(n108), .ZN(n19) );
  LVT_CLKNHSV4 U29 ( .I(n45), .ZN(n67) );
  LVT_MAOI22HSV4 U30 ( .A1(t_i_2_out[28]), .A2(n108), .B1(n39), .B2(n108), 
        .ZN(n38) );
  LVT_NAND2HSV4 U31 ( .A1(t_i_2_out[3]), .A2(n108), .ZN(n63) );
  LVT_CLKNAND2HSV8 U32 ( .A1(n52), .A2(n51), .ZN(to_7[1]) );
  LVT_NAND2HSV4 U33 ( .A1(t_i_2_out[1]), .A2(n108), .ZN(n52) );
  LVT_CLKNHSV6 U34 ( .I(to_7[16]), .ZN(n24) );
  LVT_INHSV10 U68 ( .I(n22), .ZN(n23) );
  LVT_CLKNHSV4 U70 ( .I(to_7[11]), .ZN(n22) );
  LVT_NAND2HSV2 U81 ( .A1(n18), .A2(n19), .ZN(to_7[11]) );
  LVT_CLKNAND2HSV3 U82 ( .A1(n14), .A2(n15), .ZN(to_7[22]) );
  LVT_NAND2HSV4 U83 ( .A1(n58), .A2(n59), .ZN(to_7[5]) );
  LVT_NAND2HSV4 U84 ( .A1(t_i_2_out[5]), .A2(n108), .ZN(n59) );
  LVT_INHSV6 U85 ( .I(n38), .ZN(n73) );
  LVT_MAOI22HSV4 U86 ( .A1(n110), .A2(n108), .B1(n36), .B2(n108), .ZN(n35) );
  LVT_CLKNAND2HSV8 U87 ( .A1(n60), .A2(n61), .ZN(to_7[15]) );
  LVT_NAND2HSV4 U88 ( .A1(t_i_2_out[15]), .A2(n108), .ZN(n61) );
  LVT_CLKNAND2HSV8 U89 ( .A1(n63), .A2(n62), .ZN(to_7[3]) );
  LVT_INHSV8 U90 ( .I(n35), .ZN(n76) );
  LVT_CLKNAND2HSV4 U91 ( .A1(t_i_2_out[25]), .A2(n108), .ZN(n50) );
  LVT_NAND2HSV8 U92 ( .A1(n50), .A2(n49), .ZN(to_7[25]) );
  LVT_CLKNAND2HSV3 U93 ( .A1(t_i_2_out[21]), .A2(n108), .ZN(n84) );
  LVT_NAND2HSV4 U94 ( .A1(t_i_2_out[24]), .A2(n108), .ZN(n54) );
  LVT_CLKNHSV2 U95 ( .I(l_ctr), .ZN(n106) );
  LVT_INHSV6 U96 ( .I(to_7[20]), .ZN(n26) );
  LVT_CLKNAND2HSV3 U97 ( .A1(n16), .A2(n17), .ZN(to_7[6]) );
  LVT_NAND2HSV0 U98 ( .A1(ti_7[22]), .A2(n111), .ZN(n14) );
  LVT_NAND2HSV4 U99 ( .A1(t_i_2_out[22]), .A2(n108), .ZN(n15) );
  LVT_INHSV16SR U100 ( .I(n30), .ZN(n31) );
  LVT_INHSV5 U101 ( .I(l_g[31]), .ZN(n30) );
  LVT_INHSV6SR U102 ( .I(to_7[6]), .ZN(n28) );
  LVT_MAOI22HSV4 U103 ( .A1(t_i_2_out[9]), .A2(n108), .B1(n48), .B2(n108), 
        .ZN(n47) );
  LVT_INHSV2 U104 ( .I(ti_7[9]), .ZN(n48) );
  LVT_CLKNHSV4 U105 ( .I(n95), .ZN(n94) );
  LVT_INHSV4 U106 ( .I(n69), .ZN(n79) );
  LVT_NAND2HSV0 U107 ( .A1(ti_7[6]), .A2(n111), .ZN(n16) );
  LVT_NAND2HSV0 U108 ( .A1(ti_7[11]), .A2(n111), .ZN(n18) );
  LVT_CLKNAND2HSV8 U109 ( .A1(n91), .A2(n92), .ZN(to_1) );
  LVT_INHSV8SR U110 ( .I(mux_bq[31]), .ZN(n20) );
  LVT_CLKNHSV16 U111 ( .I(n20), .ZN(n21) );
  LVT_AO22HSV4 U112 ( .A1(ti_7[4]), .A2(n111), .B1(t_i_2_out[4]), .B2(n108), 
        .Z(n32) );
  LVT_INHSV2 U113 ( .I(l_t_i_1_in_0), .ZN(n107) );
  LVT_INHSV6 U114 ( .I(n111), .ZN(n108) );
  LVT_NAND2HSV2 U115 ( .A1(ti_7[23]), .A2(n111), .ZN(n33) );
  LVT_INHSV2 U116 ( .I(n108), .ZN(ctro) );
  LVT_INHSV2 U117 ( .I(ti_7[2]), .ZN(n36) );
  LVT_INHSV2 U118 ( .I(ti_7[27]), .ZN(n46) );
  LVT_INHSV2 U119 ( .I(ti_7[28]), .ZN(n39) );
  LVT_INHSV2 U120 ( .I(n93), .ZN(n41) );
  LVT_NAND2HSV8 U121 ( .A1(n84), .A2(n83), .ZN(to_7[21]) );
  LVT_INHSV4 U122 ( .I(n47), .ZN(n74) );
  LVT_AOI22HSV4 U123 ( .A1(ti_7[26]), .A2(n111), .B1(t_i_2_out[26]), .B2(n108), 
        .ZN(n40) );
  LVT_INHSV0SR U124 ( .I(n110), .ZN(n42) );
  LVT_INHSV2 U125 ( .I(n42), .ZN(t_i_2_out[2]) );
  LVT_AO22HSV4 U126 ( .A1(ti_7[20]), .A2(n111), .B1(t_i_2_out[20]), .B2(n108), 
        .Z(to_7[20]) );
  LVT_NAND2HSV0 U127 ( .A1(ti_7[25]), .A2(n111), .ZN(n49) );
  LVT_NAND2HSV0P5 U128 ( .A1(ti_7[1]), .A2(n111), .ZN(n51) );
  LVT_NAND2HSV0 U129 ( .A1(ti_7[24]), .A2(n111), .ZN(n53) );
  LVT_NAND2HSV0 U130 ( .A1(ti_7[7]), .A2(n111), .ZN(n55) );
  LVT_AOI22HSV4 U131 ( .A1(ti_7[0]), .A2(n111), .B1(t_i_2_out[0]), .B2(n108), 
        .ZN(n57) );
  LVT_NAND2HSV0 U132 ( .A1(ti_7[5]), .A2(n111), .ZN(n58) );
  LVT_NAND2HSV0 U133 ( .A1(ti_7[15]), .A2(n111), .ZN(n60) );
  LVT_NAND2HSV0 U134 ( .A1(ti_7[3]), .A2(n111), .ZN(n62) );
  LVT_AOI22HSV4 U135 ( .A1(ti_7[10]), .A2(n111), .B1(t_i_2_out[10]), .B2(n108), 
        .ZN(n64) );
  LVT_AOI22HSV4 U136 ( .A1(ti_7[8]), .A2(n111), .B1(t_i_2_out[8]), .B2(n108), 
        .ZN(n65) );
  LVT_AOI22HSV4 U137 ( .A1(ti_7[18]), .A2(n111), .B1(t_i_2_out[18]), .B2(n108), 
        .ZN(n68) );
  LVT_AOI22HSV4 U138 ( .A1(ti_7[17]), .A2(n111), .B1(t_i_2_out[17]), .B2(n108), 
        .ZN(n69) );
  LVT_AOI22HSV4 U139 ( .A1(ti_7[13]), .A2(n111), .B1(t_i_2_out[13]), .B2(n108), 
        .ZN(n70) );
  LVT_AOI22HSV4 U140 ( .A1(ti_7[29]), .A2(n111), .B1(t_i_2_out[29]), .B2(n108), 
        .ZN(n71) );
  LVT_NAND2HSV0 U141 ( .A1(ti_7[21]), .A2(n111), .ZN(n83) );
  LVT_NAND2HSV0 U142 ( .A1(ti_7[30]), .A2(n111), .ZN(n85) );
  LVT_INHSV0SR U143 ( .I(n109), .ZN(n87) );
  LVT_INHSV2 U144 ( .I(n87), .ZN(t_i_2_out[16]) );
  LVT_AO22HSV4 U145 ( .A1(ti_7[19]), .A2(n111), .B1(t_i_2_out[19]), .B2(n108), 
        .Z(to_7[19]) );
  LVT_AND2HSV0RD U146 ( .A1(ti_7[14]), .A2(n111), .Z(n89) );
  LVT_AO22HSV4 U147 ( .A1(ti_7[16]), .A2(n111), .B1(n109), .B2(n108), .Z(
        to_7[16]) );
  LVT_INHSV2 U148 ( .I(rstn), .ZN(n95) );
endmodule


module regist_1bit_24 ( clk, rstn, in, out );
  input clk, rstn, in;
  output out;


  LVT_DRNQHSV1 out_reg ( .D(in), .CK(clk), .RDN(rstn), .Q(out) );
endmodule


module top ( clk, rstn, ctr, a_in, g_in, b_in, po, ctro );
  input [31:0] a_in;
  input [31:0] g_in;
  input [31:0] b_in;
  output [31:0] po;
  input clk, rstn, ctr;
  output ctro;
  wire   po1, ctro1, po2, ctro2, po3, ctro3, po4, ctro4, po5, ctro5, po6, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n1, n2, n3, n4, n5, n6, n7,
         n31;
  wire   [31:0] ao1;
  wire   [31:0] go1;
  wire   [31:0] bo1;
  wire   [30:0] poh1;
  wire   [30:0] pov1;
  wire   [31:0] ao2;
  wire   [31:0] go2;
  wire   [31:0] bo2;
  wire   [30:0] poh2;
  wire   [30:0] pov2;
  wire   [31:0] ao3;
  wire   [31:0] go3;
  wire   [31:0] bo3;
  wire   [30:0] poh3;
  wire   [30:0] pov3;
  wire   [31:0] ao4;
  wire   [31:0] go4;
  wire   [31:0] bo4;
  wire   [30:0] poh4;
  wire   [30:0] pov4;
  wire   [31:0] ao5;
  wire   [31:0] go5;
  wire   [31:0] bo5;
  wire   [30:0] poh5;
  wire   [30:0] pov5;
  wire   [30:0] poh6;
  wire   [30:0] pov6;

  PE_5 pe0 ( .clk(clk), .rstn(rstn), .ctr(ctr), .a_in(a_in), .g_in(g_in), 
        .b_in(b_in), .t_i_1_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .t_i_1_in_0(1'b0), .t_i_2_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .a_out(ao1), .g_out(go1), .b_out(bo1), .t_i_1_out(poh1), .t_i_2_out(pov1), 
        .t_i_1_out_0(po1), .ctro(ctro1) );
  PE_4 pe1 ( .clk(clk), .rstn(rstn), .ctr(ctro1), .a_in(ao1), .g_in(go1), 
        .b_in(bo1), .t_i_1_in(poh1), .t_i_1_in_0(po1), .t_i_2_in(pov1), 
        .a_out(ao2), .g_out(go2), .b_out(bo2), .t_i_1_out(poh2), .t_i_2_out(
        pov2), .t_i_1_out_0(po2), .ctro(ctro2) );
  PE_3 pe2 ( .clk(clk), .rstn(rstn), .ctr(ctro2), .a_in(ao2), .g_in(go2), 
        .b_in(bo2), .t_i_1_in(poh2), .t_i_1_in_0(po2), .t_i_2_in(pov2), 
        .a_out(ao3), .g_out(go3), .b_out(bo3), .t_i_1_out(poh3), .t_i_2_out(
        pov3), .t_i_1_out_0(po3), .ctro(ctro3) );
  PE_2 pe3 ( .clk(clk), .rstn(rstn), .ctr(ctro3), .a_in(ao3), .g_in(go3), 
        .b_in(bo3), .t_i_1_in(poh3), .t_i_1_in_0(po3), .t_i_2_in(pov3), 
        .a_out(ao4), .g_out(go4), .b_out(bo4), .t_i_1_out(poh4), .t_i_2_out(
        pov4), .t_i_1_out_0(po4), .ctro(ctro4) );
  PE_1 pe4 ( .clk(clk), .rstn(rstn), .ctr(ctro4), .a_in(ao4), .g_in(go4), 
        .b_in(bo4), .t_i_1_in(poh4), .t_i_1_in_0(po4), .t_i_2_in(pov4), 
        .a_out(ao5), .g_out(go5), .b_out(bo5), .t_i_1_out(poh5), .t_i_2_out(
        pov5), .t_i_1_out_0(po5), .ctro(ctro5) );
  PE_0 pe5 ( .clk(clk), .rstn(rstn), .ctr(ctro5), .a_in(ao5), .g_in(go5), 
        .b_in(bo5), .t_i_1_in(poh5), .t_i_1_in_0(po5), .t_i_2_in(pov5), 
        .a_out(), .g_out(), .b_out(), .t_i_1_out(poh6), .t_i_2_out(pov6), 
        .t_i_1_out_0(po6), .ctro(ctro) );
  regist_1bit_24 pe6 ( .clk(clk), .rstn(rstn), .in(po6), .out(po[31]) );
  LVT_XOR2HSV0 U2 ( .A1(poh6[0]), .A2(n30), .Z(po[0]) );
  LVT_XOR2HSV0 U3 ( .A1(poh6[1]), .A2(n29), .Z(po[1]) );
  LVT_XOR2HSV0 U4 ( .A1(poh6[2]), .A2(n28), .Z(po[2]) );
  LVT_XOR2HSV0 U5 ( .A1(poh6[3]), .A2(n27), .Z(po[3]) );
  LVT_XOR2HSV0 U6 ( .A1(poh6[4]), .A2(n26), .Z(po[4]) );
  LVT_XOR2HSV0 U7 ( .A1(poh6[5]), .A2(n25), .Z(po[5]) );
  LVT_XOR2HSV0 U8 ( .A1(poh6[6]), .A2(n24), .Z(po[6]) );
  LVT_XOR2HSV0 U9 ( .A1(poh6[7]), .A2(n23), .Z(po[7]) );
  LVT_XOR2HSV0 U10 ( .A1(poh6[8]), .A2(n22), .Z(po[8]) );
  LVT_XOR2HSV0 U11 ( .A1(poh6[9]), .A2(n21), .Z(po[9]) );
  LVT_XOR2HSV0 U12 ( .A1(poh6[10]), .A2(n20), .Z(po[10]) );
  LVT_XOR2HSV0 U13 ( .A1(poh6[11]), .A2(n19), .Z(po[11]) );
  LVT_XOR2HSV0 U14 ( .A1(poh6[12]), .A2(n18), .Z(po[12]) );
  LVT_XOR2HSV0 U15 ( .A1(poh6[13]), .A2(n17), .Z(po[13]) );
  LVT_XOR2HSV0 U16 ( .A1(poh6[14]), .A2(n16), .Z(po[14]) );
  LVT_XOR2HSV0 U17 ( .A1(poh6[15]), .A2(n15), .Z(po[15]) );
  LVT_XOR2HSV0 U18 ( .A1(poh6[16]), .A2(n14), .Z(po[16]) );
  LVT_XOR2HSV0 U19 ( .A1(poh6[17]), .A2(n13), .Z(po[17]) );
  LVT_XOR2HSV0 U20 ( .A1(poh6[18]), .A2(n12), .Z(po[18]) );
  LVT_XOR2HSV0 U21 ( .A1(poh6[19]), .A2(n11), .Z(po[19]) );
  LVT_XOR2HSV0 U22 ( .A1(poh6[20]), .A2(n10), .Z(po[20]) );
  LVT_AND2HSV0RD U23 ( .A1(pov6[0]), .A2(ctro), .Z(n30) );
  LVT_AND2HSV0RD U24 ( .A1(pov6[1]), .A2(ctro), .Z(n29) );
  LVT_AND2HSV0RD U25 ( .A1(pov6[2]), .A2(ctro), .Z(n28) );
  LVT_AND2HSV0RD U26 ( .A1(pov6[3]), .A2(ctro), .Z(n27) );
  LVT_AND2HSV0RD U27 ( .A1(pov6[4]), .A2(ctro), .Z(n26) );
  LVT_AND2HSV0RD U28 ( .A1(pov6[5]), .A2(ctro), .Z(n25) );
  LVT_AND2HSV0RD U29 ( .A1(pov6[6]), .A2(ctro), .Z(n24) );
  LVT_AND2HSV0RD U30 ( .A1(pov6[7]), .A2(ctro), .Z(n23) );
  LVT_AND2HSV0RD U31 ( .A1(pov6[8]), .A2(ctro), .Z(n22) );
  LVT_AND2HSV0RD U32 ( .A1(pov6[9]), .A2(ctro), .Z(n21) );
  LVT_AND2HSV0RD U33 ( .A1(pov6[10]), .A2(ctro), .Z(n20) );
  LVT_AND2HSV0RD U34 ( .A1(pov6[11]), .A2(ctro), .Z(n19) );
  LVT_AND2HSV0RD U35 ( .A1(pov6[12]), .A2(ctro), .Z(n18) );
  LVT_AND2HSV0RD U36 ( .A1(pov6[13]), .A2(ctro), .Z(n17) );
  LVT_AND2HSV0RD U37 ( .A1(pov6[14]), .A2(ctro), .Z(n16) );
  LVT_AND2HSV0RD U38 ( .A1(pov6[15]), .A2(ctro), .Z(n15) );
  LVT_AND2HSV0RD U39 ( .A1(pov6[16]), .A2(ctro), .Z(n14) );
  LVT_AND2HSV0RD U40 ( .A1(pov6[17]), .A2(ctro), .Z(n13) );
  LVT_AND2HSV0RD U41 ( .A1(pov6[18]), .A2(ctro), .Z(n12) );
  LVT_AND2HSV0RD U42 ( .A1(pov6[19]), .A2(ctro), .Z(n11) );
  LVT_AND2HSV0RD U43 ( .A1(pov6[20]), .A2(ctro), .Z(n10) );
  LVT_XOR2HSV0 U44 ( .A1(poh6[21]), .A2(n9), .Z(po[21]) );
  LVT_AND2HSV0RD U45 ( .A1(pov6[21]), .A2(ctro), .Z(n9) );
  LVT_XOR2HSV0 U46 ( .A1(poh6[22]), .A2(n8), .Z(po[22]) );
  LVT_AND2HSV0RD U47 ( .A1(pov6[22]), .A2(ctro), .Z(n8) );
  LVT_XNOR2HSV1 U48 ( .A1(poh6[23]), .A2(n1), .ZN(po[23]) );
  LVT_NAND2HSV0 U49 ( .A1(pov6[23]), .A2(ctro), .ZN(n1) );
  LVT_XNOR2HSV1 U50 ( .A1(poh6[24]), .A2(n2), .ZN(po[24]) );
  LVT_NAND2HSV0 U51 ( .A1(pov6[24]), .A2(ctro), .ZN(n2) );
  LVT_XNOR2HSV1 U52 ( .A1(poh6[25]), .A2(n3), .ZN(po[25]) );
  LVT_NAND2HSV0 U53 ( .A1(pov6[25]), .A2(ctro), .ZN(n3) );
  LVT_XNOR2HSV1 U54 ( .A1(poh6[26]), .A2(n4), .ZN(po[26]) );
  LVT_NAND2HSV0 U55 ( .A1(pov6[26]), .A2(ctro), .ZN(n4) );
  LVT_XNOR2HSV1 U56 ( .A1(poh6[27]), .A2(n5), .ZN(po[27]) );
  LVT_NAND2HSV0 U57 ( .A1(pov6[27]), .A2(ctro), .ZN(n5) );
  LVT_XNOR2HSV1 U58 ( .A1(poh6[28]), .A2(n6), .ZN(po[28]) );
  LVT_NAND2HSV0 U59 ( .A1(pov6[28]), .A2(ctro), .ZN(n6) );
  LVT_XNOR2HSV1 U60 ( .A1(poh6[29]), .A2(n7), .ZN(po[29]) );
  LVT_NAND2HSV0 U61 ( .A1(pov6[29]), .A2(ctro), .ZN(n7) );
  LVT_XNOR2HSV1 U62 ( .A1(poh6[30]), .A2(n31), .ZN(po[30]) );
  LVT_NAND2HSV0 U63 ( .A1(pov6[30]), .A2(ctro), .ZN(n31) );
endmodule

